PK   �PkT'��~�  q9     cirkitFile.json՚�o�6���B{�I}�om�}Y�e�bC�-��H�,%-����Q��ZN��l�X�}���t�u��֔٪�Mvk�}Q���$��:�ӏG�$�e�T��Z�6����ͷ�	W�ͮ*M�dj)�V�	�$"�:Z�˕�C���K�LS&2̮�W�͜���\��#�yL3Oh�)�\��bG��s֌1�G	s�PFL��Y1t�Gi��^3���Ђ���Љ�y 2D�H=g��qJ�8�P+5'Rω����Dt���,9��[�SijI���*=�j[|?6J�j[��F)������/y�½x^�H/^"/^b/^/^R/^��<��^�������� V��7~?������b�Q|!߿�O5�O�~(�~�0�C1�C1�)�c{�����6��21��9"�М��jsR�����؜нp/^�/ҋ�ȋ�؋�ċ�ԋ�:O�����~�? ������a�1������{��~(�~(�~(�~(�~(�?�xtsB��SjF7'/�9)�צ{n���`&&�]Q�}����3ۻTun�`vMy�N�Ջ	�Y8�0S��J�XRQ�����B����\� ������c�1zdҐ5]�mQ�)���z1m�S�0q�B��D{A��D��h��}J�WT~� R	tKv�G]���ÀH��(P!*�@������IRHE�\8���S9���ɩ`r*��0G�#�Վ��qW��ŀY��xpS��CX�{l"Ɯ3�m��@�M�-�[l7|؛�M��SDM@U@]@e@m@u@}@@���F�-8Zp��9��ј��1T�U�펷4nֽ0��%�j�~�kGĥ֐қ4���!.��zi���a���M�S1<�NC�E����m���Η����n]e�b���ǫ�eVa�&:��4m��0�!���iۈ�?����mͺ�����ţr��n��{7tYW;S7�qW�ͮ�<}6�}S�g{ ����(��z��7!^0mY����Tw���i0[���X��ԟ�}�ܚ�Xm�n�
�.)�=7�l�zմ�������Cos��ۢy��[��GB�
���E�^ʽ�T%q��Oe<���nW�s���A��:^��PD�kq�z��\�����Z��r�ٌ�����GV�U��(hwvhUԫ���y,�F�0��T|��Bz��O7.U ��ӏ�^_��2�J�,n�>��w����^ � � �g ǉ!JzAnn	������E+%;IzHg""q09�΂|�� �,��J�O�S0g�#8����D�������!��3g���9���̩�g��	���Ƈ4t�Cz��!m}D�H�_8X��U��E���{ S6�zH-F||g���BE�����om��d�Z�8rs>�8&�k�T1����\�P�I
mL�m>���t�5h��uT��D�8u�����a	x��2w4�o4���z9w����|ʢTa�٠gS�e�cS|ޠ��өPR`������ޱkի���o���i�o�
s�>�ś��<pO���l~x�`L�]7�E�!w�W�wΙ)�g]�����Z�]������ޮ*��R7��~>�ص|\_���]s{�]��ұ��,kӇ&N+z���=���<^�%S���)-{#�^���θ�>�[���{��'��F�F���#֖3���˵ly��/y��S���"��@v�C����3�@r�@�����׽�Zx{=��r�N�!c���q:��;��PK
   �PkT'��~�  q9                   cirkitFile.jsonPK      =       