PK   �ZITR��j  �M    cirkitFile.json�M��Hr���!_��~Hb���ۀ��4�>�݂k��*��.�ߝAVO�T�s�	��g��2_=
��|If���y�s����}�s~�z\}��n��������O�����cwy��t�}����w�{q�뷾؟��q��t�?�O��/ꪩ���b�n�E�[��ݱ�w�.ta���׻�]A�
�3�U!t�������`U]mf�*��13XB�63XB�13XB�53XBך�
�F��Y"R ��^+�^,���^.���^0���^2���^4���^6���^8���^:����^;���^;��8Ѵ���^;���^;���^;���^;���^;���^;���^;���k�Y"R�k�Y"R�k�Y"R 6�^;+{�4KD
{�4KD
{�4KD
{�4KD
{�4KD
{�4K����N�D���N�D���N�D���N�D� .r�kgm��f�Ha��f�Ha��f�Ha��f�Ha��f��5��i����i����i����i����i���-"{�l��,)��,)��,)��,���v�%"��v�%"��v&ߞ~���yw���)������|�k��L�=�2�	K',]��h섍J',]�J6v%;�NX��Ul�*6v(��t�C����ءt���s6v;�NX�x�gc�fc��	K��;�NX��m��m�ءt�҅�ecײ�C鄥ӧ�c�Y�|���p�hwA��_l0v,��|�)?�e�|��ӯp�`���	̧������'0�>q�v,��|��4?�u�|��S�p�`���	̧ϧ����'0�>Y_`���'0��	����O`>]� Ǐ��A���G	���,��|����?X>��t�?��|��8~��`����Fp�`���	̧+��������O�x����'0��N�Ҁ��'0�������O`>]��,��|��������?*�T��`�����p�`���	̧+_�������O������'0��6����O`>]'��,��|��_��O`>]���,��|����?X>��� ?��|�i'8~�Jz��?j�԰�`����p�`���	̧}/�������O;v����'0������O`>��Ư���'0��w����O`>�L��,��|�S��?X>���?��|�i#8~�jsz�9�?�4��`����Qp�`���	̧]��������O�u����'0�vc㷆��'0��H����O&���O?}{z�/]h$�ki�c�Gžl��t���X��TV���zel]ְua�d�o*�ͩ��~_ԡ?��/v�,�m|�ͺ>�v[�<�=K�쏝s_�6�c/����fN��y4s�ǖ���?��̜��Ig���53�l���6ִ3�ݰ������8�0,w�1��M�r�39�+w�1��ͨr�[k���&[7��7�_�]R�|c�%[e����������������������O:�E\��E(��/a���W�e)hMac'���7f�#���<�r]6ߘ}W�������t�|k5�ߕ#�����r]6ߘ�#h�=_�|c�%[���7�_�]�|c�%[���7�_��Z�|c�%[���7�_��X�|c�%[y�η�E�/��*w�1��ͦr��/��)�4ܘɦJ����ld�;�jc���l��;>��})u��e/����C���u!Myl�RB�+v�����u��]������y����^�>1�h��a�gu��	%�M2D�PP��ABA/&0D�P��$��C	���ABA/�0D�P��3$��C	��*T"��͕m�nV�)�0\A����-X��p�b��`�R
�I�	��qJ)WN!&���X���p�b�ο�p���X���pub��x��qJ)W�!&���X���p� b��x��qJ)w5 ;���
��R�@Lܕ�R
V�+��SJa��1au���8��;dV�+��SJa��1au���8��;�V�k��SJa�3
1q�Ĺ��X��:N)��0Ą����R�^CLX��:N)��.;t���V�)�0< 1au���8��� &��&w{��V�)�0<�1au���8��+�1&����:N)�Jc�	��k���)�/�� W�����*.����0W���*.�����W���*.����HW���*.��w���c�-&���σ\����Vqa��(.q�ؖ��������c�.\�������c/\�������cc/\������3�>���q�Њ�>��['��d�||��/�q^.��C�Ϛ����}�Њ�>3�[�B+>���Ol}\��������81Z�յ>��qc.��C�kJ|b���\hŇV�����Ǖ�Њ�������\hŇV�*���Ǘ�Њ�����1�[b>����e��/s�Z]�[_�B+>����'�>�̅V|huM�Ol}|������J����2Z��5�>���e.��C�k]}b���\hŇV���<����\hŇV����Ǘ�Њ�������/s�Z]�[���W��e��/�||������|����2Z��>���e.��C��|b���\hŇV{>���Ǘ�Њ�������/s�Z�����Ǘ�Њ��񉭏/s�Z��[_�B+>����'�>�̅V|h�G�Ol�V�9-%��e��/�}|����j� ����2Z���G>���e.��C�=�|b���\hŇV{Q���Ǘ�Њ���r�m���\hŇV{����Ǘ�Њ��8󉭏/s�Z���[_�B+>��s�'�>�̅V|h�w�Ol��|8����e��/k||����j/C����2Z�՞�>���e.��C��%}b���\hŇV{d��v���\hŇV{}���Ǘ���4�1�Ǘ�}|��L�~����ͩ��~_ԡ?��/v�,�m|�ͺ>�v۹}�3Ufz�f��t��T��㝩2�y;Se�Wv��Lw�L��~ԙ*3�3Ufz>�f��L��������ۧ5W�I��Pse���s4W�I⹝=s���s�g��0Exn��\&����̕a�xn��7��Hh��Ǧ�'}���-��
�Zio���̚E*7�f��͜Y�r3e��̘E*�[��E*L��,z�TnּeY%/��s۵��0�{�ȽL����G�e2L�>r/�a����{�T��,�}�^&�d��#�2&��#���ƹ2L�m"�+�d��V��2L�m��+�d�ܶ��2L�m�+�d����2L�mT�+�3Y<��g���s�d��0Y<�e��`�xn��\&��vV̕����s[�����u_J]�wE�K(���Pl7u]HS۲�8q�Z�"��Y�� �]�����ү>���rN����y��/�9H(�!���p!���p=!���pm!���p�!���p�	!���p�
!���p-!���p]!���x��)�\���6V�+ܔR/E2LX��xSJa�H�0a�[�N)���-Ä�p��8���V�K��SJa���0q���	8V�K��SJa���0au���8��{V�K��SJa��0au���8���4���x��qJ)�w�&�J
w)��V�)�0�(c��:^au�R
�-<�	��V�)�0�\d��:^cu�R
�mO�	��5V�)�0ސe��k��Eq���X���xߙa��x��qJ)�w�&���X���x���������R�"`��:�`u�R
��ww��������R�`��:�`u�R�5�V��X��t�7Ƅ��5V����o'�h�q�5�*.�����7 �
�ՃU\XC���U��z��k�^m�*WVqa���%�I�6$���σ\⚴hC"��*.���%�I{6$�����7�
�ՃU\XC��e�U��z��k蒞l�*WVqa�g�}����r�Z}��'�N���v��.�1^��\hŇV�5�����r�Z}f�'�>̅V|h������0Z��5>��qb.��C�k1|b���\hŇVה���Ǒ�Њ���񉭏+s�Z]��sc�Ǘ�Њ��U򉭏/s�Z]s�[�;bN��||Y���J_�B+>���'�>�̅V|hu-�Ol}|�����D����2Z�յ�>���e.��C�kD}b���\hŇV׺���Ǘ�Њ����y0�Ǘ�Њ��=����/s�Z]C�[_�B+>���'�NO+:=����*_V��2Z�յ�>���e.��C�=|b���\hŇV{%���Ǘ�Њ��|����/s�Z�]�[_�B+>�ڃ�%���/s�Z�%�[_�B+>���'�>�̅V|h���Ol}|����j���:�$sZJ���j_V��2Z�՞A>���e.��C���|b���\hŇV{8���Ǘ�Њ���򉭏/s�Z����Ǘ�Њ��󉭏/s�Z�q�[_�B+>�ګ�'�>�̅V|h��Ol}|����j�<��:u�pj����_���2Z��^�>���e.��C�=}b���\hŇV{K���Ǘ�Њ���t���Ǘ�Њ���􉭏/s�Z�Y�[_�B+�h߶�nNm��������O�}�+OeQn�km������Ü�2ӛ6Se��l��L�L���ۙ*3��3Uf�[g�����T�� ��2��97��e�wn��\&�V͕a2xn�\&��	͕a�xn3�\�3Y<�Ke���s{A��0Y<���Lh$�ki�c�Ǔ��l��t���X��TV����܋Tnf�"��I�H�f�,R��2�Tnf�"��	�H�ɗ�Eo��͚�,��e����{�������d��}�^&����#�2&�o���@5����G�e2L�>r/�a�:r�mo�+�d��&¹2L�m՛+�d�܆��2L�m;�+�d��殹2L�m��+�d��F��2�1��s;x��0Y<�Of���s�Q�&���|̕a�xng�\��1Y<��`���,^����~W����>n�vSׅ4�-K	!�o_X��>k~�����Kwxzx:w�ǿ�>���/��������o�����������)zO���$�V������!�E�;��<HQ�r_��)~�Ί"�P^8`Q������OO?�o�x���D�8����d���wɉ�������IVM����r���=_v�>�:�Ɨ�.O���q���ۋ�o����{ϟ��Y"��Ha��U\#�Y"W��f�0\E6R�%�p�Ha��Ul#�Y"W��f�0\E7R�%�p�Ha��U|k�"�'Q>��)@�k��F����Q�Fo�X9�:*@!�k��f����S�FoY9�zZ�Ԯ�RV�|�8!�i	�S�F�Y9�zZ�ԮƻzV���@=�k�񾢕��%PO�a��i��@=��zj��U+��	���
��v�0��r ���]#�7��@=��zj��-r+POk���5�x�������v�0>&`� ��M�zZ�Ԯ�'�@=��zj��V���@=�k��i��}��6@=�k��y+PO���5��ċ���E܆�i�S�Fڱr ���]C;+ @=]�Ԯ�+�����z�j䯲O�8pz�2x���|�.����!�c��]ҍ��C���	�����ď��/�8~I�;��e���p��Vv����	����%�����/tIg:N��'0_��s�?�O`��%�8=$~,��|��"}M;�PhB}ƒ�!�BpB�����N&�P�m�cH��PhB}.��!�H`B�	��b:��+�	�&�����&�P��cH��PhB}��!�P`B�	�z:��K�	�&����մO�	�&Եti�
M��.��wL�[&�O)i�R�>&�P׻�1�}
L(4��աcH��PhB]gDǐ�)0�Є�F��!�S`B�	u}Cڧ��B��4:��O�	�&�uu�!�O�	�&�5�ti�
M����>&�P�b�1ğ���}JE����)0�Є���!�S`B�	u�.Cڧ��B��c:��O�	�&�u�ti�
M�k���>&�P׫�1�i�
M�k���>&�P��1�}
L(4��8�cH��PhB��@�_��/E�}JM����)0�Є���!�S`B�	��Cڧ��Bj?:��O�	�&�^*ti�
M�}`�6�O�	�&�6ti�
M��w��>&�P{�1�}
L(4��=�cH��PhB��D�_5�/��}JC����)0�Є�+��!�S`B�	��Cڧ��Bj�2:��O�	�&��jp״O�	�&��쎉!�S`�t�ϫ���ڶ|�F�ڶ��B��g�t@����8?�8�9?鼚9?阚9?�t�9?�P�9?�,�9?��9?�䙛?��f�	��J7S���d�}Y��5+��r�y�nѕ[����n��+`���6T��LL7~��fb��R�~�W�`��+Y�h��$X4�J,�%�mzo���q
�)gM�+ui��+eiY:��њ�馥�֔�v�\&`M�k�e�<�v�\&`��k�e��h��k�e�L�v�\&`�D�2�D0W����}��LL7���fb�5]��5���r���n��+`��tó\k&�[��
�O����ƕ+`��t��\k&�;N�v[31��)W����J�f�b��t�\�+���K����({	E}���i�c[�����}]4̂_�Vo���婋�ϫ��WK\���^RS�V�?U�S�?M���6��6�iu�0PG�+:Xt��p��Dg�:��uF�3J�Q�Rgē��w�%�G@����ΨtF�3�GgT:���ΨtF�3*�Q�Zg�:�ށΨuF�3j�Q�Zg4:����htF3�i���f���y�ט5/c�<�͕.�R?��[���[��J�'3x�^�w�ޅ�����=����F6�����?�����W�_���C�n�����S�p�|>�%��+��>���t��}�O�ݧ�/\o���t��^�����v�]|��Ï�����?_�������Q��V����|������O�w������Ë����~;^�#�*���~������ϧ��s�ܟ�x�|���ٹ�ߗ�s\}���?��v�/����r���^���7�9�N���?�����s�;�SE�oO������/�~
eUo�z���h���kN�m���!*���=�O�MQ5��q�$~��ݩ�}��m�߭����e�xx���0r�z�o���V/�����C���~���S�>�wu��,��_�j3�����Q�nG-�F��:\U�����^Ӫ6�a�v�J_M[b"?�m��Ճ�\篪A�ن��2h��������0�����/��r;�m��f��ګ1+�AkS��He=�l�op:Xe9�l�W�r!y�	�+7������4���izX�OK�gz\������~S��%_��ao_��ߧ5`b�סt����./���?��籪ȧ�I���#D�'y�/�����n���ws'Շ����!b�V�/�b����&���P��8Ѷeu�b�?"��/8D�����6����M~T�~�7oŤ��(g�a�jc�j7U����T�e[o�t����7�7���z�a[��M�[��}�>֯$�[�l�0�p3��æ^tbX�?m�c)�M�%�whӣ&߀��J-���wR7#��Ǐ�J�������7�N�q��!6�&�ζ}=���$�ԸI�t�$]:l�n<�m������q�t�I�t�$�xxݮ_�D;Sg��Mҥ�&��a�t�A}[��?��K�M�%�&ђQ�d[�/ζ~WHd<��6n�v���)��~=I�ۯ'I������o��w{�`b�I:l�(5IV�g�m�ÝM���&ɒa�dɨI���ĺ�Z�'�M�%�&ɒQ�d�ȿ~=��,6I��$KF�d�9�3�R>m박߷x�/M���V�������b�9���������Xl˾,u_ǯm�?�w*��B��S1��E�#mxK����7������PK   �ZITHy"F4 � /   images/6e5c9ab7-aeef-495d-82e2-c4e48423bc54.png4[4����QB�MQb����g�j�l��c�Q��6�U�ګ�J�{����{�YR��|���s��ܼ���g<'����}r���  ��|� ����� �I�g��P�罹~�ϯ������� 8���_ZY4�$/�d[�/��?H�Gr~���f�w��8�KmYW�zn�� �RU�h,����s��7���k��Hv��yl��/e�ϻי��6�E��g���X�J�p"APT%��"��113�5d��X�:c�(H�LyD
�>S�Y�l*/��!� WAZg��q3h���ǧ^F��� �L�[T��4A	��bE!�L�a�wۍ��)4�`����n�LO[����Gs�wF$
b�5��3xh����
>��o�h�NQ,ͭn�l[�nL�E����t�N٤�B&
�V�0@ �O?�_���j�G�+�\W'�6��026�I��}�g8�p�h�k]�����,8���詧7��GA�#�Q�* �p�k4���Y%R�%&&�d,¤<2�Ihii	ܛ755=S�L�a:��H�ʎ)�RLMɪ�V�aIHȤg]Hp��^Ng�Bl���}_o!f�>����r3\ϒ��)�����P>������	1����	��:AI�3w�v0e� lp,Q����ޞ�L&�4Ņ�)--�=� �o�K@����ˆ�:���t�x�� �G�Ɲ�I�(jݗ��ɹ�Դ����搾&���&���S�5Z˪(/O���M�F�F�>������\X�+q�8č*3�Rń�L������GR��mQom���EP �_%7�h���&����)��� �cYN���i�J�mt�LX+���V=��T�m��T�b(�L�-.��Ss���֨��5��T%���|-�\VsL��!R���%,,�O������B�z}RR_r=Ju�|i�5���"%�E�wwqV"��S���ʓ���50��U����8����~��C�bi~�u���)�?�H�Fc9Z�t�餻���qC.aMN3��2�AKS�J���)Ϻ҉/kr'{ZI�������о��w ���R6�I�����������0h�&�k������E78$���FZF�TLX  ��t��>�k�M�8�x��L�~�����wb�w�8��D��}CU�͈CW����n\2d2u`%kro�\��qF�$𿛜}���t�1\U���~dA|Bg�i}u��o�O�����p��C�@7&��Z3,4�&^|�
�{�U;Ɋpw��A~]3k* W��q*	@��Lh��ߢ0���E����I�\q3?<mv@�V=����{�8�x*� ����؞�P ���dsٜ0�l"�F���[ 1���wǻ��#�Sf�.���&3��؉r����6�`�L4m�����c�Q>�:�$	����m�Y�f�hj7�I_�_knQ�v#SO�e��RD_v7����^�"D�h��LO͹?��`����ϟ�hR:�J��=��G�ܰ�<}�F�@�����	��ɿ_��Ձŀ`I�'a4���$��ƕ*��C�����=v���3"Lq�~�ި�4t�����o[�����֦����!����qؒO'�bJgL:aM�N��w8��YH��P� Ff����`�Q_ ����u����A�s�l֘��IЊ{�7���0q�3��ss�{G�@j9�oπ�de7�r�7�%456� $E Q�L��l����;;��q�mQ��ُ�1�S`�:cM����)���ܜ���\?�t�Q�<�=0عn�DP$�gȒ$�>*����600 |=VRRr�4V�,�&e�}u��.���:��HZ�,^bbj�<R�>6�����_1
ĺ��9t@���	r�1ɋ�01��Ff�^�����;��w~�2�B�f� �R���Py0�XH��If��E!L��KzI�O�3d�T-��@?�OWG���\��D����Q�� 瀤 ��w7��4 %���x�_�O�	ydJs�x�������O����o�H��$�g��r7j~��w�\���������ȳ$�7�0����~���?�~�����LJX ��T������ �o97ݙ�O�u �h�������}�̰i�>�dw.md3--�7;�5O�Q����z�\�Y����V�"9�_&\��b
� 4<a�e�)�e�b(�@�a�����A�ѹ]�G0�%��}��7�w4��-.�#F0�،m�(�l�����
q�J���x������O�T��z���F��Օj���Z��|�ͭ�~5 i����GMp%-9`餩�鉆� flll�q�Q
D�!D4�1kr$��DꃣH���J�9��ɓhD�I�j̰""D�W�`q)�$عޕ�1@�@���@MDqv���i�|]���Mz�w �1S����Q��I�#��'4(�.Ȼ�/!�l���x�_g&�t3am�)���`Q��ɣ	JY��$�?�U���y{���cɌhnltő$��kIER�>U�k8[Q��$Ƅ
|�e�n����c���3�Z�-$x����k��F[� xvb�{��ү���\��?�VsA:P1!{�x��R[QF�> �s���j0�6����r�ؑb\����dv��m�ɣ��Y2��c.�c(pF,�]�CJfX)����v��<�g�6�{8�"��Ց7Q'�;{��4���;��o f�?\��"!JՏ{s�t=��U`��K}��"�G������ �����T����  �aJ����f�Uz�ĲI~���A�n����,\�O�i�t=to?&��$l@nQ���jf�a�ƝYT*B�C�p��+�B�#���CC����w�XX*�������5^bP�����@8U����hE�����#�޽ Kc،���䤑��n�J�J���v��"m ��G��r���|����*F��aʲ�$�wu����2EP>-"#Dr|�	��gg$OL���wgqn$���\�p��"~������Lߝ"R�)�Ep�O0����B��s��tHy.��c'�F����tuu��v��#�0�v�>�덞���pSVq���#�d�_� ��[�qLOu�qug&n` nr� ��#�Y���RH:u�����%Y*2gX�z,�
h�I����s��'���dT=�I����� ��	`�\s?d�]�)�0�G�V/b�ѳt��ֿ҄�7 3;��	d�~�7�������1��yo`0�+56�̝2\�<R�x��KC����O�
���0�����+R�'�54��.&��K�`�&��cv~t;����T�Dq!O��:��*�Jw$3x4����N�|��$��`h��)�g�����s�
`3: ��|�y��4��PB� �I����� R> ]��>ȇ���[h�ߵB9�.�a���7,h3-d"<��򆆛�7��3A��3���O-��3Z^"�ʢ��ӽFeC���	ă_�D�C�>�^�0��Ȍ�!7�˸ܟ�iF6�nHڀQ�t�Q�|Y��:�4���I6�Y"�~7�v����p��@�w�C��,��`.j ���� h�5��&l�����z�9��Աo7�5���|8�'�H�|��]�z�[�y*^QÊ;�:�{W�u�o>(����=�����2@c�M_����4U��������(��I�!�Q��)��& t�l���n������$�a2t?] ?a�z�wlD�j�]���ͩQ,A'tes�A��{��/O�c��X{�vv T��fzpB��ߕh�����Z]���G��G��ߧB9����;��o�<!��}2�	N?E�~5)�����^~W'8�@�E�ۮXQ#�Ȼ��*�Шʎ��0�q
333�=U124�}�ɉ�f��7i���%{�	�R7�o�A��ֺ}������'{-Oޫ������zމ��E��p��˗Է%�?����o&A���dE�~�����i���E��kMC�j-���j!�?9_ Zl�\��Uer��g���~"
�I3��l�����պ'�oWi"�8������Q)^��Ϲ�YI��<db8B��q�MA2x��������N�9�64�6	S���H:r.�H���L^��j���Gy���Br�l�kW��??�(��e�����g�W%_��l�����;��L�nܺ�|���e�bb�s�W�y��V�����Sn��Ѭ��q��������f�!ޡ+�O��с���?�{}�:lq׍�-/wV�_�GY��Q��%O)l�t ��~��H��a��:���-Az�s*��d�P��wA>���[/Tg�Yr�K@�RY��V�+���jo���_�����,��½�II�b�m��=M�V�P$�󴷰����s�I�my�y|zݠ�ɍ
2� S�/������]h@��9�{��yC��7"
���T�*�o3'��$��#�>IF����\���&����~�>;�"�?��/�%��B���a��	�F�/-� ��ƍ�D�-hkw��qyԦ�r���{��ԞeS~����z$ć^�б����	s�ƶq�Ő�J�`eG�)o�sx��X�9b��Kö�,^�	�_�3�z����WH~�?%��|�J)$"�v,���5*�à#�TNȱ�?G�K�m�w�qv��Hm{�x�Z�����i�ܰ�R���;8�"p"�!���^����V���Y�B���A��ѵ��Ty�����Ds�V��6�ٛO���O2�ӕ,S+7 Xܚ�Y0��1��˞;���f���t�N���-ߟO,T����y�:h�dz��7����A�	Ēl,�c�����hjj��_ݳ�f83���,=�3lʽ_g�]C�%c���$u����A�	I0)8k���}+��z:��:����ĸ#<��X)�KaŠ=��Z��V<~�v�B�Zy�*��\�$��*��`rQ���zN�/�>�`��Ľ����GG��$]���<��ϵ�.�u$�΂4ޮA���v�xn�<���g��+@����RP^F1���u�Q̟/�'v����������XAx����e�d�����P����Q���D=�8�j�\W���9�~,�HT�~�EQ�F��7�QL��{��#���n5s�� �U�ܩ�"��~�S!�j��w�y�A���d�ɜ��g�P���
o��w���9��_q���:8��0^�kx���[J��E�0�w3��^�1*F�3<|k�sƷA��ȣ|�-A�/	�f	���R��Ж��m�91���Ŭq-��j�7��ho(Tuy����3���{b�h�	�� W+_czg�l&G��'vF��`m�8Hs��< #U"�~(�p,M=�CՖ�xV���F��������N������i�������j�Uq�m�B7gGdA���Sqۜ%��gj���AK��j�@���\�@\��E�R�I��4��6��^��ƌ��o�~��0���l�77�P?\Z��TX�F�S7�.7��w��U&u�|@'���BNq8|/Gs��01 �o ��:=�����+�d�NPmv����=��:�7���`�E�|��_�58��_��L�g�}�|�+��kd ���Q>a�W�[�غ��0@��S�@�4O��$���-��#H���f���Gvw�}F�F��<Rm�Q��X�����)DB�k�ɞ\��E����8fp�����o�e�~�aWPQ�$�4YVL�<��#&��"b1�2y�|��q3���Un���??�+�\5�sC�O
��+�\L�\D��]P�l�/���tɘIR�zT }G����M��Cff��t:���r��@��~<�\�C�d�ae���?�a�kr�us>�s���u)�݀���a�F����,��/)��̶�s �lƟ��V�3�jVQG�;��䡬��n�)��e���	Vi#�]��#e�\_w�"�8���Vr���;5EiMM���v�2�6I"edE��Ý�m�m�>�/%�aT��m>�2�RRN�}2��f��~�K�/�guk�|�\�&to����	y�Cŏ��(M�b��ʄ�͓������1��Ѹ���	�IWFb�0�+�lc����Ӡ�Yd"���j�ιx�Uw\o����Cg�-�^��D�1�Y\�HW��@��N�� � ��K m�5�J� l$��V�tJ}Ԑ��,q�B��FQ�Rz�m�m�P��}��� �w���xâҬ��}�3|�� DR��H�}"Yw�~�SK���EЋݍ�G,��Ծ�6(}6��Y==��Xc����SP ���8��r�ؗN��:��|�Ʋ�B>U��h�R_B�G3�,]-��{���4�E�\V!>�nNs)2�z<����}��p�{�6���j�������[V�{p�RqU����O���Lu�[{���0��m�2o핖�xP0p
�I���!P8.�MY�=���W��fުT��Sr��
���[ j:83�a12�b���s���d��j�@r:E��޴~y�1�r2C���?�����t�ʥL7ɔ��N��U�sm��g�U�___h���y��h j���Y|[k��]?��{)�i�e�=s�����H�<|��d��-��_hjneqD�YN u�F^�Č[7V:u�����]�$��ۧ��^(܍��݁���9�$I6I��g,����/s�q	k` �ˇ},&&F�.��$%%�u?[�4��%�ӏ����2J��?i#����������Ο��h��ҧZ^~����o��x�΋%���%����y��Qo�~Z_r$s,\~ז�B�m�|��e���O��k�f���lo�8���o1�@j�SE�wZ��5�H��YKd�h6@�?$�a�;��m?����9�}̶�hJ�;��`��1_W}�i���'t������ψ�i(x��ȩʐ������0ea�f2�,R"��u?�C5ض�L��6S�������2AO��|�����Xq�Y)�R3�e��n3�,o ����^��_C���	J׍���ꈠ��[W޿����E���xDw�_��w�e�*�e�Cf���ϕ��7`؝���g�#�Vs�	��i�z�N���C�i�o�.(I5|ԏp?by��3���O��*<���|xV�_U�(9��_�~��ϟ�q�E�˄X������3�k\���AP*2�?��'��ƥVR�����^����FTs����3=��Y�!� Gʸ�PpmJ����OS���[Nw��M���?d����9.�/�"��⇂V~$=1t�ݟ���כ` D�'ґ��-g<����=m���2f�tq`|u��tq1�{y0�+y��n�=A*��/���"1�k� *����2��H�ԓ �������c'����,�������{�AOX��N���9�)%pI��-�@��*����"W��E0�����z1�N����6N�͑-�1�
������ܴ�i��b�P��GǺ:a�n�J5W�%���N�~�V���ڤ�I�e��n�u��_?{Ɯ��*��Swu��C�����}�o~O�9�5�p&�Y�� .�� 	��/��*8f�-�맬��W	����N�z���jXɋ5[�!�*A'�����7wZT۾VU�@
_��o]�P���n��|��em���nyqA�(�j
ttČYu͸H?�����VD}m��^vS�ESx��R����_S<.�W)0���"A��F%.��A���)��#�G�x$�֔��(x�ݟ0Ձ��S����*�'{�X�sok��2�Z�����Q�������O8:mQ��@�)���W�D��9�ީE��B� ndi�n��Ȕ�e(�x��$�!upck�n�i���bHz��@�E�;���^2*���f���]�!�PX�C:z̍1$�����kTJ�5XC�g�����Ԫr��$��������+�Svml����7[nٔ���G�#{�Պ&��$$��M�[|uYə���P�>J����ܝ��Y4��Ʒ��4\`��u_eee���F�����Xx_�x+��h"3�)�H�+:�������&����G�v]88&���Y_yy���N�Yg��K��*��ZBZ���)���c�R��M#I��M74�X��ܣ��5wZ
ۏ��Ƚ����2�ZgZ�4�[�n&@\g��R�ݶl���'�ě���OU#.�ތ֬�=�ܿ�����]o�ذ(Tn�ozy�ro���H��^��՛��O �t��Du�(�/���|]�~�U/���☋�݆�0�u��rĩ��l�'�SSV|��,��\0(��>/9O(���/mh�6ˡB�"*zE��������-Y����C1�3�ي�K�-��>� ����N0�Cm��˙8���p�ĭ��̫uհ���=sZn����:CVrMťn�����������1����~�l� x�����bEA���@�e��)a�os[��GK0�;�70��������U��Q_���J:N ��|�l�������EnS���Uo`����_W���t�2�ņ��Յ��W�Tr_NT�X[}v뽍�R�	;8u��qoٜ���~��a���q�]wu6�T>T1R��`-x9�W6��E�c��[6�Ygk��D?i�-us�۟;�0ܛ�?:�im��n�X��̝x]F_�#����{�Y�ٍu��'EL�D�B��P��v��"ǌ�u�������GB|�e����Yz/�gE�����Tnֿ��S��^C
Kf0l����o���o�.�eT����g�a�W�/A����'x,_��ʹV	�v�x�.v�C���h��ֆ?C��#��)��`Ii��U��W�S���ٷ����|��
A�2cUr���3t�V�E ���ه���3�Q��G���g���r1��kЇ�>p� �8�k��K�\�D CEMM�K�RD�m�׶�@���#����\��r_V0�KD�\2�l�x`pA�H�D(X�!]�h�d-���L��g����T�����گ� U���r�ҋݩr�dj�Vdta��=��Fdm�?�s'�Ď"�;������M8=g�l6	PȎc�a�_�}ϡP�/����N8-�vww��4*����O�����yfz� S�W��i����,\�ϛkFYgq�+wâk�ǣnX�ZZ���EK �p�m&"���Q2<&�
	5�*r�
B�i��^��	�Y �`^�}�=�{/Ocb^����\m犇�[P���'<��Һ~��]X����Y��l�Ƥ����>�H���4�{����ؠzΡ��`���&�2j�,�ᵘsDH�h��09q/bc��˄	��M�M؋��f�*�j�|Or����5��,"��̜��wH��h������6A!@E�G��
��Ww�T|�*�}ow��w[v[��g�4�����6o���"�ۯ�� �3Y!N(L3���-A�N�^�eW�U���k�eB� $c4�qmc|�׿I�7w�|��g��?Xll,�B�'�o�r�4��ؿZP��y{߿~m��ǯG<M��U^'��}���r�@u�ȃϏ��)����A�5#�%����u���O���<���XT4�~ZRqkVks��Rt�*@'#�����?ށb�WkW�mk�rb�C@��&`�199��$a��&6����7�w�@)Łd��vqƂܹ���_�m_������^��V0�hE��$t����JcN�����\��1�3S����
��cTz:�U숸�\R�	y� Y"|���|�w���ʳ�x�w����u�-Mu��3����j����R���m�
:��xE�̍u9YdO������'�o)����oN���6�� ~����Tm[�s����������5���t-�)E�Ul#�D�^����V�_�����#>$ΰ��˝���j'/:]���֍��	�B>�沯���[�� ��ɜuL�Ֆd���Կ�p��Z2	<
��:*�36^-��8��������r�^���,�VV�ݨ�t��{�x��N^蒑~Sy�7��.������>Ì"�X����E�%?2}�\��������q�ǒ�U��ܑ��1���� �^(p�����F3Y��S��Ͱ��2s��X5�w����[<0_d }]�w����B"5ͤ�W�z=>�3N�.��(�����3�d{{{w7K�����mȺ����� �[�}����1��:�9$.>f���l�ʼb���!������)��zpd)�K&�4մev��e������/�����>�:�jJl���x�� �B�b񖪪��Do�$$�:�|�F�:�+����8ѯAD<m�_���>��G�v�e�Y�o�MU,6�ګ��~~�Q�d������{�/�7FQ�ڋ��Ks�k�_|�T�t�-<�mz:�6� ?Ra�X5W��
��֔OK45n0���c톩���/��X[�%I{p�ԗOJjVe�O�Z�50��v�v
��y�٠ �JNv���rs��R^0��!�)9�x���h`���8"��`�+9��z��7�Sq9�W����ݭ������Y��%��:E�
^X��z麻��p����ޮ`g1kD.�0�a�I\j�D+�X�^lu��^CŴ;���_o��K�Y5���31�/ݝ�>��/X�h��Ɉ�)��[�?t�Q�q�	L�$T�0H�ՠ*�Tٜ�X�4��\��q;� ��<�gbf�mmU��Q2Xp�v[j�O!
A�|�0~L���`��c�(�z��T�ݖb�i	����աxRD�����13������VP�G���u�I�W���6g��z�݂s�#܈�w������5�l&$��)�H�L��E����bYFf�8��Ip7t��M��鱣A�[GqoC����{��¨�ў�_0�2�(g�q�s�w�IN�|�UB�%��~�9�)���,f�j�S}�ǡTS/)�[ cq:keK3���dJ�u3}��%������J�����(H��Wl�#���b����d���5x�;�G�� ���UP���k���y(�R��>�p�J~e�Љ�<������-����μvD[|�ڵ|<)@�v��N/pң��P�^
��L��? vl��E�I�h�z�q��6� 	�[�~R�Զ�WI����d���3��w'M�v<�5?� %�l*f능=��xC~m�r8�<f�x�Z��9�Dg����!R�`!f,t'�#b&��������Jk�O�G̭,�7n�U��{��|�Ql2]���	�5>7@��J�I�,�-心�]��:	{`>^ɤV ���Xj��F�a��zUѐb-����$bT�䴓��?���Rb��HU�b�?F��z<&�����擨��x@������&Z�)��DXxPT:�nK��%
��w�2��nz��6��ܤJ��a�ơ����gD_4��Ew��WH�[�ȋ��1����o�R�&^�(g����x�]���� ʧ�I����>���a�d�k�F�׼o��~���8���m��48��ݡy`Sʍ�OH�/������*���{7$^�!� �A�	�'�*��o���/�G��	��
`�Zw����\p�*yҝ����_�Sԝ��Er��bƟdg0���M�����^�ڣ�����踺�T؏���>O$s�	��v�����-����}���FA��-�Yi	��?׆����0A����Fp���YH,L��R�Z�Z��{�V{
�N6Ze�M$¶�nRu&S�hZ� ���VHh��5`�Eis����6[��^VM[����?~�="㝏d�ی=ut���n�7JY,��2���	+���¼FGҤgZ����9w��nz+�R��gt�ؗOXF� ed1�W �O���{�7�X|�Շ�J{��D�BEfd� �[�:�A�ëm���/��}��������Mej&ɓsi�܆�4���-в�r�8i��E\�Zl��422�1nCA����Y��OJP�|�/FĈ���-5��A����z������ܜ�����q��6 [��.�ן˅���v����X��=/őW�o������D�|�u�H��P"�]� ����U�4��OF�3v�u��C�k6si��G&�6X0���6#��s�NN�tuS�1�5��;�Ź����.��G$n:���=�\���3������$�36V�G��M���<L�k����ڟ��
w���9�䤤����d6p#Q�����F�5�7Y��*�H؁Fچ�l�>��^��h�px-dfX,�3�!�!$Dv��h�ǉ+�o�`�#�^���ʩ5n�J�E5Si��+��TAB4��7x�oOI=���D"뤞��"�B���6I	��6�bH��Gp!M��(|L���&v$�|��P��k��^�^y��Ē'�2�g�r[��>����ZNSZ�YKX���jMtA[VD|��(mB�"sh�Aŏ��y3 +e�#������ B[�����vB�mH~lrj���Mmo�(�(�G>�zw[�agvJ��Ȋ�:�Z���5���ZcfF��x�v�w��%h<ü:݁��G~3����#Fޏ	l��<o�O���*�P	��]����ќ}o�o6���������J�i�S����I�9��۳��c��������o����'���b������hðH��1�[(ou�3��׷�	Jt���w6��;�T1Y̌��'��͊�����I|MI�s�zG}t�%靤�E��\�o�α�[���HJ�u�,?�28�Y��3���]�cT�0+6f��'y'�_B��Ĺ@��������p�����5i�Mh������S]�7�j����&f.;Y	�Z����$��4dX)�>?�����,�;�_�7c$�y]Rrr�O����R��㎘4�4�u��E�a�����8�B,���5al����*z�)C��?��u�!!�S#�BHb�1��J��͍�B4�[?K�T�c���9��
�q���n�����6�������_����y��wP6U���k1���n��0>F�˔=Fm�7�E` 3�[M�x��2򢌴o����T�,�����r	�TT(���Xđq������bw���v`���P��i��+�K�w^�jhh������B��qy�&��0�����	���O�N�'�W�֗��w$�0����0���#��>37�����kZ�4�|}�]B��"�cӖ�x]�s�z�	0tK�勲�H"��5��`>�N����xW�gaܐ%|�,/�V�x4PF7g+8&-�K�W�Ov� {`(r�����u��p��5%�⛰��J_(	�u�OsK�x���Ʒ��q*t�%TMР�G2�����u�B+���0��i�: ����t%���M~�ee�0�͛�N�-����[�h��X�1��1���nl�o*�s��r۶���eg�6jU��������*�2r]q��.��b<H<]<�D�'=B7��U6�x^�s̥�GI��(ڱ�ŕ�%,������:,�N��n�`E����Q��R�p�����)�2�/��^��"Z�|�n����M���MZqf�7<� ��W �OT�q����TX��xd�]�sh��d�\V�ߧVO��[��0�1�	tj�t��H0��.K�@���[z�<̲0�k�X��-T?�v#��d���[rA� ����ӯ4�I�a h��)��z�/c!4\֛�y�жX��~��]9�餦���>�wz�#�E�,�W7o'�Ҵ��12 ��]7U�
�:�s/�f��m���(MP�2�T������W�u�ߙ�071�RTI�S�����$�,��-�l�rk+��y[�W6�w��
ٺ�W��g�z?�e=�"�z�����p[���c#�������k+Oĭ��"v����)��$OK�ڻd��&x��
��D)`g���h�ij%)�꼌K�˫��$[�z���jt���c������]��{Hp�
9m��
����fp���M�i��#���W�\�r(�">�q��G'',)�-���]��sc�6���m2$����
���hĮ��}�G��h��W�{`&TF�v�ַZ��4�+v�y�u�-TH�)��<q�k~��~V�3[�$�~JQl\{�s�p��|��Eow9:����}*l��-���Izt߮�Mm3�4�`1��=�^��	���œ�=���Q�:���n��y�?jݑ��a�N�M�o�*�$%p�fM�|��▍��U�x��7�h)��̦���X[��>���*3��� 1�b8qwN���n�2	:�-�7.ˇ�<�<�<�����O��m��;򽐼VG= �W>"Z�֞��ü��2"�2��|��2��U�eS�jaڗf��-��u�'��;��Qh�T"�y�J���4loB�ڳ�����})���˅'��B����_3\�r�Y����kOW�Ԏ���J���ss��g��t)���!1�o�rCw¹$�k�.&q
��4XN���W��mA~�+�.��J'��S�-?�u�C�^��n�N_�/���,����W�ӝ��n*��~(#oZŃZ%]�ժ��:�	>��X2I[�]�{?�����<�:�1�l>�<��yoW�	��'��zU���G��;]�?��1�3�I�T���D��ݪ�o1rm�n-�{�l�Ν�o
%�^�s���HJnh�=������;���B���{�V�bq���J#6��&��	�f֪�7�`�+�U/��z�u�m�������9_�{�N��3��X�/�Ü���~xN�h��i�q���#��M�ֵ8�%B��y�J"[R�a��T�`s����^vP�� ��{l���"bbnؓ������=�=�aM���Com?W~���L}9���2���o{�a/����`2L��A\\��ҿ?KW�[o/��ݻ�hX�u�*������� �h
��ʹW:��#���:qU����˞4��X}<5<n��x^�Z��M}�-�h��/Ith�-��� �fc�כ|O��Q/��͖d<�m�?��y%�$tt�e���f�(���W\m���01Xx�̢x�5��w�6�Y�*���T�M��u�@�JA��G.�����~���ǧI݄fN�0I���_U;�Ȱ�KЙVL�[Z>�H����z�
��)µ��
�*�
YW��jK����l"��Q��Tn7�mz��y�'�Lea�YDĿ�sW-7	nG���{����hsCn�[2�Q�&����
hr��]O��Æ�Չ�y��Ё�GE:���3I7��ˣ("=���ة�G?�ώ���?�9ɍ��wU���]��}�a�½�w�s�1�I<$�z���mooc�J�~�hZ0*��>BA��we���$�`�v���%c�:@��ԠO&r�����_`Ʒ�o�?,���"�*�z��?P�������+�}�7rw�YZ�/�s���,22
�GT`!L��bch阛��t���S�?��=s'�z�W�e�^�*	�]N?�Ň�M7�I��%1З{��0s�~��ҩ��y\�C^r<����ks�b��`G�=m��Kƪ���%'L�H�4��6m���mC������ܫ��W�d���&����;l�G�]��E� \�2�#W��|�MMb���R����?$ ����e��	���G�$��4�ۉ!�V����3���i	�G����g_,;&�-�ܺ��_�#~\��Eق��!�r".O���@EcgC��8v��Cþ���1[j�Aq��r����;��#d(���j2�q�[u�ʟg����ho��n����"
Wkɦ�'�h�_�]��r,:�0���5�	:��~�zV�%�� ����Cd�+���۷�s��|�wr�$b$/�#��9r���l}P�\��F�#�l^e�?t,�����q�?T�63�zaFRp�{��י����K���=���]]ܶ&7���{U�8.-|�1
��
1�7�pS��F��}�߿�7����ޏ+���:����������,'�8�!-�~�)ť�������P�Y�Xy��e|8p-ƤM�ϒ��Z_�g|��u�HJKW�af�n\�ֹڵ��l�8���{���[b*?��e�c�}|�D�D��m���簕f�T+��#�G�N����4��_���3��O�n�|ka>���='qu�@����Z[�o�UAE�j�0��#��l�)B�F�-��0�hld4*�>�DʔM�g�y����fM�'�����Y��,C�J����K���xS��P{ꢩ����N�>���Bc;�I�����d���#�2篯��rY�܀h,�/���j������A������k����2)FH�tw��
�&F�t��F���%�@āĨ��#"0�c�t�o~^���Y��m�}�s�u]�s?�4��0�w�dge}$����� ��)��`O�4��*�,�V8�竪�F+�$��V�"f�Ģ������啘i�c5
z�h/�w�d����'4l�翅3󄪠h�wP�0�^��{�?l3�SL�&ךd��'E�}	�hx\�O�od�|���++��'e��d.��~�p�J��������"�ήF�Ppvs��	�m�ݙ)��4Ξ����g�悅r8��/W{�C/G\w4�/'�V�,:�N>����1�}���*��J'v�:���H��W�Ѧ��!���s���p�^�y����|����oi����!J�.U�����H����B1����+���Ë����TW�_���mǨS7a4>������'��zOE`�z����6�wZ� ���n��,/{j�N���_��Jg�I
�������tSH<�5�d���̌��k7�6��B��/�n��{72�R;�w#8���^kr<�����N	��R��p8&�����6&��V?Z��j�Eھ9Z���qldK�";
�j��U���ͷ��N�Qf%~A&k���!�+(�O�x���.��Fv�5�'ُK��3�E7`ڳy��߯a��G�!g��n$ћ/Ȟ~��f:��N�Uaǽle�G�_�[���׋�����W���q� �hݴ�����yP�/�[H��o�D����w�Rz7c�ao�����N"��kS�.��7&��n�aѰ��Ӕ��������f��?NO�f����,β�j&-\�(��Ϊ�n�<�p������¢���˥T�,��I!3��ſ��GG"�/V�E� w=d�Z4��>�PL���o���)Y���C/@��qt"���,G��ŵ}���l�Y>9ZʖWgԽƔS��u�A���Ȳ��,��
�|�C	R���y/�~彏��&�W{�����FX��i��	�wݳa��Qo������gês������j��53����W�2�ǡj����+�BH��pR�����v�5�"�@��	���UGo����k����v��UGؾo����Ѡ�sW!�qcξ_+++��0X燜s������'(:;_IU8��(��Hz��?�cZ�;�RAj1ԉ?�+�z��s��f�"�8Gggg7�_-�8�J��OVo�8�����2Ҵ7y��t�Ej��0�=vFs��_^���Z[{{�����X{��"%�n�q�D@f~Q&�1����BE�,�84GhM�8��p�l��������^�2z��p�ޥ�M�� ��?�;�a��9�u�L8 �34:�O���e��z ���w֥�Ɉ���z�|a��T��ͷS�}E�}�ĳ���ݯ�D���C<~L��_�s�([>ٓA�Qݛ<����γ	� >�d�5<
Zf/h�{���CƠ�G�F��\���M�O�ĄO�[����΀�k͎:I�pD�K�ceG��_�֛š�]�3��1�A!!��O�����j"L�������[��K,������p����WE�A��ޗ�jg���{��I�jRHl��qp�_6
/X�p~�I5%�!�U�W��)�1ػY��?����GC$��Y�7c�)M���Ư+������U�k�8�W�>�����2�O ;�y���zE�QD�6�3������a'dύj�����䳗-w߼
+M�=�['��:e3�����C�ݨ#�N��4�X�1�'��P�I����AW]x���H��;�;��e|6~Y�L�\���e��ݙ�*�Ě����陼�WOhp��]5�M��-g�����y��Q�u7a��h�y�WA�:��渢���E��y�5�ww�|�J�)��^Z֮5�b�����Sӈ�jW���l1Y �����wӣ�S;O$�n��G�BOxR��-__�m	K7�%?N\�8~�}B����[;ܟ<�n�o�y�o@��~9y{]�p���>�Y��M��E�����͒|�=-66��aV��B�����H��Jh��Y}La6��S��-#��eإM,�hWt��c^�̲S��$"%u�Y���p���ŭ�3���{Wq���n��:j��E�j~]]lg�R�xv��:�H:�Ȟ��a�!z ��[�m�F+�S���=�U�ϓ��$D����&ws!�:�X���Ϛ����x>N��RݯXZ�=���[h�u�+/8r����秳�ۙ>AԄ����0ݝ�J�N�㎒��A�Ћ�*�:ؙ����JI�bz��ݼ�y�=�y�pJ�[�m`��ќ�Y��:!S�2ZVH�<�:vwcy���(�t*�1�Oʭ��w����NJ�Ld��ߓ?���g�0Q�����:@53�k?���">�e�[S�}Z�qI���H\�2���N|��k4����z;=Q�9�y�΋��F�~����9:�l/Pβb�qU�3N��y�H���#�;SE�2<��#�Jj�o�K�7P_����YdNT�z�����SC�_V3z^&���vi�'�,�r�h�a���	Q�V<�p�`�I���)F�t�o���������7���J��h[��$�C��r�h2MS�������՟�GѲ?��u�����+j���1��g��XYmYOj�����IK�MQ]r�쒗�R�m;�n��D���+��(�\�tl⡖����0� �I-d�	��y�$��d""���b�z�,��+�ʻf���D�/���^3�K�Q7�(1G4��'k7�3�zx�T��+����q̍���ըE`o�\����q�Q����i�3W���M�9lT�,&��NH���B֨��C.�,A�9�����Jv��3CCC��++e�����y����K��}�&\k~��ÚG�B�v�-�g����"E��w�4�h���"�!o��}=�dl\|��u���֒�a���d����6~q}�<�r���F,��6�c5��L!.Tj�����Kـ�.|�>�Zi�16U�4�La�7u(;��F+�~k,�mx�p���jZ��%s�ݗV�����k�1r/Q!y�{w7K���=kYU愽{�IM��n�{ɼ#�q6,PDi�
�^���-�m���)�N#76�=��MH7a�lw[��ac�5�������5��#r/W��ŎGx"1�Z��;C����RM���D��Blll�]R4��:�%�dX�����,~�{����冪��Ș���̖뇑ԭm�m��z����w߆�QE[o|��lUTT⚛��+v�WHY��;��h�Hц�tV��+������-�k	=J���'b�W�n�ϛe��p�W[]��,�����{�����Z�a���o��.w�'kBy1�G�����MMM�&����F�C��v7ӷ돰F����4�� 9>5%OJcY�j�����=�P��I�
� (�lr��h�܃�#�=3���+�"�����+��~s��Cb��n�m� h�0��ц�
��Qg}�pjU��q�ts�S�P�v���a��~�3"���g��R��[���unx��<�<a���sY8�p;_܎�N�xP�O�H���򞾦��R�=B�03ӄ���������nw�H�����`���5fUfwI�Mb���b����0��4e�zQ����CN�-ۮ�������Ia3U1��x��T����^�Y�We����'��Ӂ��<wK#L�-y��U��s���+��b�X3I��u���Q�R�'O^�'mo֞e���z\��x�K/M#À^C��upK�������7�}#�����k�1�l���)
[���C���φ)��hm*fXJ�f�S^e�t���xU�Q��'p�h.��MP�.��<��o9��ٙEl�.\b�
D?9q�f�ؔdz�����_Ѧ�҉��v�	Hq-��:M~����D��n3v�y9�z#��q0P% ug[6���駫����Kl*C�lP�1��g~�.�}�u���8�ڨb��p�f���4���mIQ�A�e�g���h���v��=��:�غ�UmCz���a����WfG?"4�����!=-l�E��&/!�6bԃ<,�75S�q��q��̓���O}��7��_�h����p���"��` �]lϓ�5.ee�������he%E:+̀JMKK���� 'g�&YE��K����#B��I����w��Qڣcg7�-���)
^�D�y2�u{�vƼɟ�����e٪��s���z{y�'�-/��p���S�-�ڹ�jr E�v��n��<0pS����!?�Zȶm1�������م{�p�}Vt����/-Y��J���-�׫f�(�nk�j��=Bx�%
3�����,l�_Y�(��q��˭*lc�...zT-�s1��5i�'�����^�`ݓ�����Yv�[��ݛ�^���w⿛��qx�N�����	������C�yr��8�~ۋٛ�����D��N�Az��$X���Ogӵ�v>,iE����#�U)�|�ո{ atH~8�`��A�?����|�qlꤷ�P��L��V�����$O������%��Ia��=���;����s�-�Y}Lx�I�⃌$/�X�� �uS�R�����r&��w�c�7C���jKG�t:��X�ao����>2Q���:ߝ�y.�6"
� $(����I�"��S8��T�5����cˍ��>�\{�%�,��gt��6b�����Vnjq��z� -�/=�Q�N��f��T1ը��؇q]�Jv:+����4h���ܮy��+�QF&0�)�	���Z"���?��f�N��,Z��������ɍ�\ �Z��W6�D��8X�\;,Q�-���AIISj�m�@玆!����#� ���p&l?~�p8�n���q�.;La>Ly*cXi@�(�n�['_�f��e���^>���!C��	AہY�_�ay�u�)jd���R��#{�c�G��Z�_La���W��"��NR�tƸ�$�tD�
a��_m2g�G��Ay�ӁA��#t����#w���Џ�,�.Oե*�D���tw�^���E�k>������UV�e/uo�^R�1�[^�-.*����PǪ�yH﹋��)���5��K�� ��54��8h��g�~I��˝_f�~�����?;���"HN��	��z�����u��Ө�%�^�vrh�i�wknڷ��2O4��za7^R®k�^�\BN�G�Ri���i��e_�u@�_�����B�8�`�Aa��U��a���R���蝙&~~���ufs�́5o*5�|	��&�P:FF?B�v��DC��:Lk��E�4*NR^ނ;�A:�zc�C���?7��1�v0-<a
r�ӗ�j�����#��|��v4��cH��@=��P�ĞHGVW��Q]�X����>�b�+���6IR��n����_j��x+rD�?*r�T�� F�:� ��K�2�3�G^%	Q���+�Q��(ex�8+]�������Kb<����0�O+�Me�.�i��yY��z� ��t��@T���)�9F�WHy�N�_�D"�Z�R����]$�='�=�j��.�4����Z7�^��нֿ�u��q^������QIzE(��e.����m�<��,���Z��B�Z�~��	Ɛ���Z�3�IF�z�Yl��/l��ݺ@n�F�$���ۃ/�0���_d�}�"Sgk�^�%�|��V���G�2/w��>��7.!��<��<i������M�9�7C����>�Ė���)���;)��dO�F����vfl�/Y��!F�i����;؀е�L?������\Ȃ�j�+��R�R�8P���.`�CN�SI���M���CҨ)�T
�]p]�K�V���n�M�Z��8�h�	J{3�2��8%�i;,k^��I�{�t�r��y����l���^�T��.�ϱy����CF��cLO�O�X �2��! ��I�##z0�L���Ǝ�:dT�L�U������ʙ��ɹ%Q�}F�ups.��sh�q=yF����^�S��ε�V������Qq�Tr���vD�{�\>D�f�L+I3}c&(e���^�S�$�z�|E��r$�҅z�/u�������yqqj���_���r�;ӈ��Mê�r.ۡ����S���
�X䕣r��͓;~�PM��v���y�	\u(�ʶ56b�OhP^fU��99�V�_��������5�N]�3Z�3��[Z<�uw�O/ܨZ���{�7�����x�{߸���p^��� /�Q�nƔ�Q/%�=6VV+�c���* �c栮�t�R~�����F?퓶��~��ˁ�Qd/}YA�������t�NR����^�ț��4�,luR���l̪6�'xfF�=��Mf��ı�<mQtL���Sw�@�'��&UKY�%�
��/�]�ك����B���&o��{�5q���Ž�
p�D}E`L1oQգڊ�Y����EL��MP���F���Y�b�G��S��&E��[B��f�!�.O��}��(�Dqd�M��1b��D�������su̗�J�
e ���.�l��%���X{�ޮW(��o���� ]&:��� s8&�+����"p�O�]�0>_�;G�{����_�~�xާrŤp~��9ޑl��=���j�5����1���\��@f�6ۋ���a&I��y�^�u��B5����:�շ�]�d[^�4�qڐd�W�F2o����'
t4����y�6�m����7MC��Q
K�Ln�/����/�l�!��ɭA1/�6�ι�����0�B� �[�[`߻��rw�����B;����ORF����R@��e�C|�3v
�Uw%),
��,J�L���> ߥ�-�}0��^3of�����<�#�a��f�.7I��*�X�z��c(�|�Q��5)��;�Xd�}���+�M���M��,���(DS���x+�@�Wݑ�g�sH�Q��)ۤ���G�W�V�,�e��>�M�}J���Cg��(��|XRR2>>nXu�+k�9Wb���N�"���ۋ�W���͇����V�bc%�J�J��ve*���n�H��	$�:���y8�Q3���BZ���}��^/�=" ��S�̰���+��	���@�P~�b�O��N�C�<ڨ)�]�XV��413�TQ`�	'c�K#Y�-������%�ōD0��"�I�.�Ə�Q�0��=%6q)�F5`TWAdp$e��\V_��K��E&�1$�
%+U�ñ&ao��,����qEX)C�;����$b�$�j<��qB��O���8�S�آ�=�9��G���{ 4װN{\�^l-�?���(^W�T���-�ɴhQ4y:D�S�����.U
���x5E���-Q=�K�^_���N����*�PE�����p/Y"��nQ�i΋=����6	/�Ǩ�����櫎��wf|��᣸��I���A���J:w���[��Ԇ�����ncRîWF����]&~�s[A%Ö_�ׯ����U�F��V�����?(*"a`�Ë́{ӊ(��#S�T&�H�gZ��Z����K��m��S@��r4�n��� ����i� 0g=,�c��x���q�.���Dzg���p��c�W��'_6@��&��ܼ0/�˸�I�9pI��I+�D�'��{�^֔����Tj���).��~W��QI_�C��F�Ʌ�Iz�KEu�`���>�{}_����֯��1F-4Y119v�φ!������,s�h��
�5�
�R�>�8q� ��gS���--����V��M�Ҧ���`�f$5�x��F�|12Y}e����gvʝ����~��ҳ0��0��pR�He��rd�:zd�@@W%[_���''p�q�}l�2~���:���)��B).����,�e�5\ ��(e?]�U���[�*$}���T�} 0T�[VD��N�f*���uH�x��ơ�C���'�<|<���{�+���x/*ΑG�`EU���$�߄�A��jd�C����h��ɷH_�>
��]��U�6�m�#�%�Q�PdW�[�7c�OXٮ/��\*��l��{�T D���J�XP&���<�ZoefuQ�6���dŘx���j�Ց�X�gQ&�|<~hVh��*�[��H((h�'�~*�f�|$�x&���t�R؜ �͠�H�D�'|��x���)I����#�B������A폏Շ�J%wDMM�rH�m��mW���}T�&�����{Ľ�R��66R������Kd9h�KX&����!u.1		z�h\��nɱ���"l�;(rdċ�s������ۼg?�9�����\^^FC�V�_n
ue"�xGM�$�Y�%�'� @Q���}��)צ�h�n!�-����H��癵���VYY�cE��E�-f~ۦU��0r����\�L��}l65Ί�k��aH�\�� H����cJ7�8uz8˯��:(��B���S����C/`1�9�ǉqFt����#��IwX10�r�E�{�cf栲�I��Un�E�R�CN��5��/��B^e|q�����0�n�yʵ���H!�â�߽*^A�Je�q@#���b]�}}/3���I���
f�_W��:��#0��K��f�Q�ɚ�j���k��w\R���T�|���H�&�P��n����k|�zq�Z_N!4a�f%+�I�,,ޏ4��,��M���s�¨h]�]��=�&� �O-,��t�lvU�>Z���W��WO�)F(
��@��#�Pw�A��8	��U�Aa�<�
-dctB����/�w�8H��a�6�4EkK��_��I����EA
~�&�hrI��~)�w���W�7�Z�uQ��.I�ɴ%�޷�𝅵�u�8:^�@ z�-�6�K��B���]���ّ�I��V�8�����!��vR�uaޗ=�+������%�h�U] �n�G���!����u��Z7��)-�3E������AvX
�z*����PIޜ ��R 0�\�D x{�DL��B
k�BpJ�*Շi���ۀ��jr.���@����9�Q��`S�.P�.�
�y�V��U<{��n&g�9bw����uKݻ�['��rٗ��+�������9u�1��d�j���z�+¤6��KV��7e��s8af��X)���;��)��՟��R>.8�k���]5�l�y�݃������N��MO���>�׷Y��+��+��^�V�{�G�|ÉP|%M^ͼ��9AZ|�̺��iZz~�0�N��'x�I�y�YM7�H�
�B?$Jѕ�'�7���n�F�좁3;�)r��LL�Kmj72bbb���[X�w��m�(��a̛�����:�`o�S,�2�<���&tp7��X��!9����{\@@e����G<[���ϲ�%Col�/C�B�u�^ɻJ*��\Y(���+B��f(���U�v� +�Qq)��Bv�ɘd��Z`Z��+~����w0O��c T����b����4��P��Ӧ�!�c%�] �
O�`�QT��T�s!q>|���:��E /�jc�1"2��Y�7VV�o!����-w�&�8���3i��Qdb/��F�?�n�" ^<���[.&���5����D�Fx�&�I�H�&�᧠�Xl��O�]�2��A%���@��î8�j�I�C~
����#�>�T��[$�-	(��$�^�F�:Oh�O�E%�j�y�cr�n.g�i�v���AҒt�ң�%�aN�a��`��AR��/U����'ť��)dB~ިF)�}�M5��Mc��}�7h�O$_EՎ E��J�8Sd��ԫ`�tUr|�K'�䴾���F+������}�l����A�E�`�(�_VV��<�����x�$%(�e�} ��"&���f����Y�G�����i�����)�34|i�98����~!׎�nEd[1U|�����v�r�7�k�����v�x���ރ [�H�G/�"ݴ�X����QOd��?1��H_ӟ�kG��t'h�����qX�ɸѿ{�M�ۦ��|����#$��0�]I��J���֟���+}�潢�y������!���42"	�������N�X*�\6�R����D� �%�˲�z����3�uNwY�A���`ET���v�?�`�O|\%��؋�g�ښ�ؖQ;Z[]�U��R]�9Q��Qk)l��`{�-�������5G,F?��3V���G_)p��^���k�H=}��&�{*�������.�����7�W�,��
�lK���KZ�"�أ[0yBZ����N�s}�0A��w�>�Rk*d��N�\��O��+E�� ��Ŏ�GK)q@���$�6q}�z�"q�
'��15�;��X����W��p$��1�d��[�%���Q�$W��h	�#�[fݛ�OԳ>eN���b��j��8'��ݦ�.ߓ;���76�6������9��E/!�:;���P�2
�D�?���T�=��J%}��pj|ҏ�E���YZ�;�/,�m�O�.9���+Y���T�I�8��rţK4�+�<���� ���BRR&�T�s��;~� gD�~�oV!��+�4v��k�*�3�h*:>�o�cL���]#j�gV��!����&J�Y�>��ws���%eĝ�@/�w�f��7ܰlf7a���q\��+nB�r���v]�s�a�t'��]�Ѓ>��'<�j�rZ?$�.;�XJ�*�șmj��3>�;�����;�d<<�fvN���@~��l�Mhh������#��
����ᧁ�kk�.;}}@��&����g�j�\�l=p�iE�4D!e���G�fĕ[�,,-�z<��g[|��q|�{___���aw!� z�����l�� ���"�^[fO���9y��xi�{���e��
g?���&	�3B������4�D�l�އ"i�H ���5�����e;B��C�y�v>���$L&�.��H��Cn6��"V�I#���Ӽ�=�XK����g��3�
+��.5�P9.�dȝ��Ҕ��̙O+ȟ�Q��͖s9x�W�;�������y﷯������&L�SqΑ0��3|��WĐ���K��	MW+����/]^w9:��p&�M��r�\V��Z�!S����W�b*�v�l@H���=�Ȭ��lA�����L{�1��8Yp�U~�����k�TY�h�}s˗0��X �#~�hJw05����C�o_���������r@��MK�u8,�7�W7��8�T&36}�]p��]���&�OuvP��vȹ1��L#ܢ���عiFUT\zBD?��l6˚�Z��M6A�X�*F9�#�gqI2K�cBI�.1q� �8?�|s��cn�ؤ{{5�͟�¢��		�,�ߏ������\���l�tl����#���W���\V����}9&3�O{��q��!S~l-�R��R����f�J�z25�+��:���1~�P�5�jXU���Ȱ�Ŷ�����g��K��.�v<��9��4��y��H�$������	G���|�m@.r�+?!Bw���Ż�����%��III��>�{�ˠ	%�md�!���D�y�>N̘����L8}��<�|�Jh��ι>s��=��]\����	9��b5����x�<��:Y����p�b��}�m8h��R�X/p���~�n)���H��wU�im,ˡ��yԓL� �����+���滞����8@J��cq�f9��v��/�G�O��p,ы�E��0��yj�&�5:ÇTj��ٵ�N+�-�mk�
X�L�^��['q�f��to����\t�|��_p�%�	2)6nS �t��IK7�}g��(�o��,9u$k�]3��2��i�4��!�r�-���ܲ�<���ێ���[=���A��,!` |}��g�"��AG����b�)�1
��99U���q�c���n|�����4159_�Qz-�t؅�3�4���$�����4Ր;[ 4��ҶXRR\����@A���@����9�дq�W�m7Y(s�0�*��i//{�h3�]3��V5ϫ^�"�8)����L�l��������6^霚P����F�oR|�d#)�bi?&���ɂ#�'��f�!�(m��g{蔙�>ՠ]�]�א��/rww;յC=�>�DO�h��t$�?�?Ϣ�H�qo�Ғ�"�*\�	1^y�L�2��z��w��/v;�u��!bZ���3�z$3���z�-�k:^xJ��ut����~�e;�W>��4j��/\{�� �吮3���/>xf�Wn_�4��v��JE�!��f�ˣ�����˟�IW��y_��Z�x^%���5���M���^u���������l�zH2�^݄v�"����@I���_R�+��ȝ����dL��nDDD$kߓB������Ϣ��l���>geg����I�������z-Kvx�%`�q��[��Da�>����?A�V|���ӯ���j�>̆�~t�e���UG"B�� �Ȓ���]���$�����B@1zT��kJ��u$|��l0���$yf(JD��ɪ ��Z���~�f�V��s��6��H~��HТ$)6ɂWW+w%g#���Ys3}�j�Z%�H�CY��b�]p��@~R���G�Y�N�c��L��İc�=��G_�Cix��C��=-���J�B���X$��ě�q�@�V ��𷓖yZO�F7ըV5���+�㺭�c�3؍�]�����9����.�ͧ���t��Y7���Z
!k;ce�ﰥ��כS�Y���l�n�
8�1�*��ZT^��]�J��ͷt�>���nll�SKDH��n�s|�AwDͻ"m��.������i�S�%��
s鈟iv�ǵ�'p?��ߢH�-L�A:E����$e>h�p&ߥ�X�Kx�1IM� >�>��u�R�h����yLj;�s��YIE��8��������uH:W��N.:��A��"�`�3ڰJhBw�:��67�j9x����#6��T�~�36�'��̝��'*zIp���JN�}Vhz��y�S�9�Μ+�K��v���L���jQ��C.X�ӗ�(�f�f%���VVK�G�&���S�؜L���z�@�+++�?��*��*�-��|�&β���3	�R{]&�3�V��,J��A���e�����U�:ձl������v��EǢI�H�:�P�0�G��2��]4���������2�j�	I�lu2t��,����p��5�����t��J[��2�,6���J��:^���vy��k�cGQ�d����355�V��A���-��H~�'�@��#;~� e���=�Q*�﵋9�V�
^S�/�tRr���c���T�[nN�����D�Nۙ�ܙ	n3zTnnn����0ŶO.//��EX	�8au�=y2����i�Ȣ	���v.�Ғ}��~^y�.��=>���VմV'�}2�fݍ���I��~�V�ܔ$�'d��V��C�a�Q�yG�:^������;�k���_3��qg���V/t�����H��\�7����5�L?��Kܘ�O	�:�<�f$��>��B��? s�b&QU�y����%
�h��lw��=8h�[$���⋈_8e����Ӏ,�\����t;xfѼ�k�{Թ��B����2l~��n��lwh�C{����Hc������nv�'1Qڷ�pL ;���a\)m-5Q�]!Y��-*���י�v���B`�n���q�p�Q�g��3����v?���`�f��f>tt<����S�3!cGj{g�\���G(�Ud|�W�Sgoo��O� v���m�])߿oR���Д�CVZ%� ��?���u��^5��]��a�պ{G��T�u*exU/gb���";Rw�6/���-�Iq�P
�j�r���p�@�w:�`l��U�F���� �����L���w���[��q�P��� �/\�Vԓ�A~o���0JQ7���⛿ɢ:n3躿�k�J�O`>~~�	��	"�����ق�޵.^8������h!�w���bL�����k�Q4����2�t�r(W�������C��������2�L�{�>�����ｻ۽����(ՀW�b�~���6��Rf%���	���g���[��kӘ �b�<<|���E&P��a#ϑ���^U\�F�R$���
���7`d���aNy�N��[xZؔ�=������,�G(��#5�MgԻ%	�Y���j-�.������Y��?��b��9�0��ղҀ.Y=�h��i�u�k F��\�DP [P��g����3��+�A�^F�O~���������z�rʒ�hv��L�	�.%��J,P �,0BT�oP3C�e��m����)���7[lգF�^/^��\�4
khl4tӎr��把�����:����e�%�9�yy����pw�����yr��	mKX�,�ƾ�e�;��=ݢ)��=~N�%�-+4��c���Y�p�(2�G.����L�������"�e�Wԛ�����Ԑ�糆Cu�+7~g=ѿt�ed�^bܚ���-@d���q>��1cc��'iXr��L�?�Al�ZZF�B]wG������/�DY� ~�U�^���d���*t#��Q�Vr��\g�}��ꐠ�ې÷�$�\�<XP��Y���X�նE��������\�lY7V�+��<��.iy:\6.U�?�\�f��y��y5P�e T2�,���^E�j��v�d�����
+o9:�Y$�W6��%��		�l�0�z�in����V�`ʊ�t!NW*(D9"��x.0lni��׬G�677�������)���l��M�	��eL�͞K�Ƚ�mj���2�kU"5*e�w�$=F�!�^^^����38�{�f����B������@�I��3�]��}z��)Ϧm��*�A��>���o&�� ��"�>�<�퐯�k�qW"mP�V��ho]�E������{�h΄?�?����]vV�N%�c�{��͟�������=	���l����{��Ml���|�*�'����<'ܛhm���r."�_���l�v11ę�Y�Ϯ�Wb�׆�B�Es�P��÷��W�2P8L�G���\2e額,��w�ש�)ܻWJ��U�_�f:�+���� _}@�������q��E�(� H�;|���2Y�(�G��&l�����	�4I�J��|�ͣ�՗.�{���h}�dd
OɌe�O%�ot��6�y������0��$�x�fۦ��}�n~�~R�Yi=#�s�ȳ�7j2�h?8y�w������;.6�����5���(�2����K�"�}NZ��=����3���ߋ@�h[E�\G�8�HYDz��d�\*rg�=��C/���&��v:V%I���5�T�52��t�V���aP�<��_�ɵMDŞ�Azec���1�E2ϋ���["g
��mu�-��@�wO��۷X�z*�|�	{zy"v��T���j��8/��p��S���,ɒ���X������T��?����m�O2q����ܧp����*`���x��9zZI�h�7��B�1�'�UbRR�-�L�ی���<�J*�nꁁ��(��o �nh�����V���^_�;��fE�N����Mo0�
���uo��	a$^`Y_��'�k/+ń�����\�D(P�J 3�
�>3�&W `����-�{a{��$h��Jp�����O�Ԡ���[|��Y�D$���
�jc�x�T_��N��!V���-o��
Eؒ�?�|��p������SC8� P�_.*�@���<�֋��;��Ii˫�&�#��4���=ҵ�e��N[3�O�݊i��5J	}��G�*}��[�mD�.:R��d�B��fɘ�gw�j,;S����5a~�I��Η�,jT�w��+6>��(VŪ(?�Jz(�juo�v�Q�.��A	C�ANJ��
	-0�9��8��M�|F�#�����P(DUb�5d�H����ZS�J)3����y�x%@��mu�ٺ�+v��Q8򸛻��!a�j��צ��w�Y47�E6QV�݄�*�{����2����[��ҡ���y�#�==��V7��t���@غ��US~O���F�5��G_7>������*����{�g�o'��M��̭���֋i��8v�x۳�I�,¾����ߨ�e���G�Ln���d����_��f�T�t4B/��fК��p;�'�v��q##�n�g7gw�����:�J���H����9���"�����4�XU>M�6�r��ͱ&Ζ��c>3���q}��t
d����f�����B�Sl��D@��1�zN��:���Qڇ�_�.�JV](HBq&���h:�h����ka	�F#���	� �Lt!z/�{�^Fe�ޢ��E�=�F��{}��;��Z��s���<�쳏�{�����,;���fh`@�W�Q0�gce��@*/%��)DO��,i?�s*�>`?���� #�B>NZ'�^u?fN�DFF�7���(���tT�a�3�c�ex�h\�B��|��S�L�Ғ5x]�>�헸Y�˲��c��]�ZQľ$'����,),ps�j,�1�S7�K?����u����!xq�a�.�T�<�ٙ��z�Q��NfeW��Dj'���8�AY�^���?��9�?�� .#)���[���ws�U�sss\��
Ѕ�Y����B3>H�F��e�,�-�g��$��Y\,���s�� tݟ�[&Y�$�Q%���tw�/�4i�ddx�����gѻ~|7�t��U����r*CxW+Ef���Jv,�����xhU�%ݼ��S�|ܧ\�?�����V�)���TQ���LS
zNj4�V�w���9��H/v0��˿����dl��|��Xa�y�m�����<uLľtn��*��}��>9��n!v�h����Q�ȉ��m����d���6�J����9�.ů�ąV���%z�ʈ���90�����,E�������k�\��#�-A�٣ߑ�Q�Ѯ�5W=��G�7y�5����d�(���2��ά��P�	�]5	{�fI���H#h�:
)�y*��(��@Wlk��̍og(ĉ|g&���x7[Mq��P������7 lex�G
,���F��ӣ���9u/�(��6�{@���,L'�H�nX�����;���ƛ��.��ˉv�����=�iB�{�UIz��?fC����۳v�\��ml$Lb�Z�+��F���@NqѼ0�rf��T��~�Ck��d�2�z;Ho1>Cl�񱤜��ԱhEpd����u@7���L�Ћt)b�!��O���eθ�#��aܦ!��XJ1u�������Q?}�-�)�CA�rP��$�%��-�8�+�E/�kȲ���:}�vV4���3�WQ���SB��,����l���E��V�&�<q����
5!��]l*
��	!�Cs���0�����Ia@�ɇ�1�1Z�O�0l6B�`"���]��������ɖ�����o3�ًj����_6��o�����u�[j*au���`t�"�~�R_���ò��w"�=�i��E��՜�͠���{���2놩���b�I����)�����e)�0=h�)غ8h�����7��i�z�i��U�����[7������Ɩ@�K��w�ʸ�nR�'qs��$0���<���;�)��y�X���Y/�oD6�T�,�uǡc(��ҁf�F���������V�������Di3XY�B��XJ��3�n&���)�E�����K}/�g�V���	"2ϐu��b�(X�T	7�Kݞ$o41�K�+�.[�s�3F.����ڧYT�2�:��C6��diY8��^8�q�}uu5�,��������dJo߲��梲XAX��ߧ�


<<<[�_��g%���NXLχf}���q�����qZT!����n��� Jwd�ciY��s��t���$i�wgy�c�3B�}!ʼ@�ҠrGWBس�_U ���I����R��F���L�h�����ѭ�f��.�~PJb����|YVLx�g�9��p)ڰ���\�_��!tY؃�ĊR�h�؏ɴ㎐ǥEE.T�~N���p�f����j7+���\v^�w�0mA�
~�nj��H4j���`�aXl�uX�{0SmG�3Q� j������o%>p���B�]�S������1??���H\������_��H�v]y�Z�e��*q�j�H y˚Ӗ��Of��
����4
�J�=��oK4�6-|�H)�x�X쟴�j�L
ۡ�_�J^Pr6�LJ�I�����n!��ي�*v}3&q�B�.Z���R��ߺ�	�&��{3>gS��^�+��u�w|��X��o�%<k�h�^����"�F19�^H�xˁK]�t%��R⁚0��3�ɸ$�4NR���<Eꗸ�������"�Ń��;e��ۓ�O�?M��'�Ҵ����&�f��&���C�E�tMW�U5/�R�}��:y{����HH���=}-�m?wj�
g���a��o��H��NqK�D��Į	j�G���D��]�x���p�✶��S�ő6o��u&G��m�	�����N*�mȭ�+�vÜ����q���0�_���=l�GL�q�����# �_�`~�,A7���!8t�Մ2�&T�K�rP�ǘ*�g�P'�z�;ي����� M�Gd�1a�Umj��!8��rA��u���;�#��U�R��8�P�uA<����W��1_��:|���KM$��N�٦C_C���#�����_Q]Sx�
_�O��1DP�dU2�WRPk^j4�~{�}�5�C��B挕����J�+�]h9[�x�=�S�". PSW'&4���5�]p~�����9m&ffIT��1i�X&���KwAZ�n������wѢN��,6����w�!K7�M+��=v�o�%J�W�r����:�{NȦLŐ�I�����<�tl�uޕ��6:�/4W6-����q<w:���~,����OB�k.�ǖ������N"_��4�r�yߎ��C�Tp�+bx�����{0LR;W�,�:���}G�+*F���g�=�B�d�	r�8��;.i�Ֆ%��(yH!py�Q�BiS���΅�t�o1�f�<Fv읮l�B�~͕���C������7�8�҂�?l����R_�eW�I�ǏFK���u�ޤפW:�s���b�N��|��";�_L�9Z�e�2�e�N��n��~B�q(1hJJ�6}�ȗ�������(D��Vj�%��p簡/o��el]yk8Ҿan8��o't^d�ݫ�tww�V���,+�����r�M6���G�����ΌM>.�)��'� �����l��?�L�N�b\#��ٟ��0]0�jA(�}|T=�.��J4Nďb��6��0p�48��ο�=�a�R�R�0�hkP<��M?h��A���'(�(g����L�k?7)�,P�B��O����7�5������䫳	�KB��'�@Vs���g7z�,���[Q(���������5e��� ��_CS���a���e��"����6�^���JP�����O��HK]M��rR_S[�����1t�q���w��Y���d�:�m��_$���D�G�.n�"O�������,��^�k�G���$�I��Sr������ԑu��N#�����l��_}�����ݵ,�/(��w���NϬq�9�OZ[���?a�Sԋ�
v�σ?�a'�sh�we�'�vٴ�A?�uC�]�(u7�b��B����%ޒf~^�pU�KD��SK�g=U��z*����TE	��?[���A��_��W�k�+���������� V���x̀��������&�NH �M�IZ�yq4;;{r��z01w�^ff��?gWډ3u�hB��,.ªIRR��#�����
I�z� ��i����.�Y���w��
�,��~-��5)���$�[��4��(Pg3I�P^�$�������<�G����`"��\ȃ��qO��
B��u�����	p���Hyh`>#D�ro��Z�؃��+`WPvƘ ���f�<I�&���~�K��
��t*Kc^G�͏�Ti��Fc��^�^��Y�E�]�<,[�D�"N���݂�O;��!
��o2�c� �dl����Qe�Z���b(���}�f�xh�W���'?�~o%�x�mq4�My��|��o*�>���5�(�ꩩ��z��&3���f����K)%|�ϔ��EXp������Q.. ?�D�<WJ%2���5���sQ�GxR�U�J���x&���W�5s{\�f(��є|� .~���g�stbM/�OG�����R������Ng���{�Rn����۬h.� ���O2�šcH��LR��P�!�wD�&6��7u*q��״�ubִgh2�4bY�I ��,k)��<�31j��`����Y��d�OQ��,U����_eQST���
��*Z�	V�h��d�Y��\�U�6},�ҢJ���w�u���+�Yb�(DMM�iwwwrr�N�H�-�[�Kxx8F�X�d��YQQ�S���<4Q�P�aic�d``����ݿ�go�/m����H@p�"Ǌ�ɕ�S0�|�K~��	�>I�k�����?���p���׭Ѣ�z��r��f�#�w�mD&>�o�F�.\(�s�Ka�!^���RsM"-�����|��?��ܚ�b}��g2W�ͦ�8a�OelO`�kR��#ąC�����yd�	��l�g)������0��y,z��@X\KSq��˜!i+ 簡��,����?���qJ�D���=������g���s����ګ<?>h$.�~駃+0��!Mȅ�
j'f�Y�u���xȋ)���3�����W��f�S1�lְ��κqb8��p�.//^h��v���4�*@�ru�3��r�7�2HS-� k�}�S�1�[\����LLl���3�e2���;�=��?��Ww�ր_���.������[m�dz'-�_Ek'�77�L`]0����W=�Kn�Y�l���z��߿���M��Ի�:sr�x�9�
ňcW��a�q9�O��y,�c߷q4��I�
���fo�mcɁ�f6T��a�ac�B��H���<�����ũ��˷�?F����3#�~ ",��ҍ9�#�M#���t�%l6c x�J�1'�<���CK܌K��M���RnZq�����"��/��F;���:��r$��:r�Q��	wOp',�2�ԑ��Ǣ��I�(�E���:�#;������k�WͶ�(4���i)[nme!�LoZqz~^��w�$5^�p���$�`^Vk�`I��T	�&1̮��@o�GY�6���z	mҭ�C^c�h�,	L�Q�p��.U���L�&o\�>?�x̢�P�;,pk��W�'Ud9�b��T	�b���`5��۹Sb�� #��bW[]mڷ��c��s�k-���%?�!P����5����% ?�����)����w�m���>J��cr%;'�^�7�א6���hT��9��<:��mCy5/˼�P&e�����P�?���`��ɸ�W!�܉?E%�S�\��s{�J�����Q_��~W�W�z�NU������{��JF�����9䖯���������̽���]�)���b�- �1�x���D���X>.��<���cKJʮ��H��l.%1�(=b�<j��,�����诰���N|�%�sWxC�͚��g�dLeUB�}�Țh�o�˓�vٳ"L",��M�?Y�SΆ��O�3�p�u�u=���qp�Jai3u���	�[�tu��y�տ� ���6-K_SR�Ϯ����&3_��7e�*llml���
vG]�xOww;
�E.  @IA��708觏4��$	�=&$.�io���yD�x*��x`��i���˶1(t�Z�I��+a����E��):��5�Hx�cQ��O�08Q��셢���F.�s&ʐ�� [���7���!�o�>�y����b�v�&�3kr��0�>\f|��#�_�+b�g�R���?'nd\�Okد�C+4�-�	�:������]�~8�s
�@�uw��{�Ľ_@���$|uvP�Q��O����9��T�]��XEh"[l>5��hGȟ��\��8�t>r;S���%y�:��'g�}ye@)�~� �눊���&��;�z�&���L�:�$��]����*�_Y�*��ƤYLb>��܈�e�6�8�P�*Y�FM���{�|�yq��q�(c�Ŷ�����5���[���#Rs�Q��_;�\�S��(D�V�9C�� ~^�'ϢEn.O���)���N�}��D��D���_$���u��$%&2�����L����z��G�F�b���-�5,������ԑ����P1a����h���1����IU�wDGK�
�՗����P�����$p������jP�C�Ɨh�̡�1��.UQ��s�Yؒ��(2�\|�S�|�P~>��Y��#c�?N9R<$)�2�6!�=�/Y�RNh<���G-���*�m��sN�؍㉁?T�(��@��YF����D&����V�p���*7��_��yMp��P4�qq�e����η�RV���Я_�߿�Y�<�q�P������{߸�G��iv4Y�)�%��6��:��i�� /}Z���#�Lc ��!�A��N�j�����',BQ�u^�����䤆ާ��=�aS�]҃�^�8ɘ��%�i�<� 2k&Hp������_�N��}B>G�,-����%$$2�6�����^g.^�����Z[[7�^�
׿6"���P�.< @�(gx�~faE�̏\(�8�=�����!�C�[���O�|�HY/4K���*V�1��M_�9�a�2���Ӿ�����:����//�s.Tg��M�7��Q9cU�T;U'��*ک�Zk���&������_1zcI���&+�*G����ۥ)k�L��^��{(F�I�������q���)�X�鞟�JS�3u�z��ȥ�څ�c�Q��݂�d�f�Q�.ss�T%��N��.m���.Q,��r�Jb����z���Q��X��(<��թ��DUI�|��3鱯_��cz���_h��QP	~D�	F���
�i�#DD���6��"�ޕ�B3��i;^e7�C� �V[���a�>��~a�<��Y	wT���-�`�k�3�n��m�����C-w��/�K\�t�����-��0���-76�A�\�y^|4/���S�ʙ�|�!7b�*d$BLH�| �o���*:�y���)����/�ŹSgEQ]]]PЃ�
ӏ�PaKx�TTPBb�0~�� )@!���2��Wެ�Cͬ��H2#X�`�������Z�A��K�9��,K|1�c뷅J���5����˗�㑡��ͫfD�Fa�5+����#���ah5S��a*��i+�7՟=�,��aur�����%������F6��F�,M��j�9�X���a��C7����S�mu�ۚxH��3�������,���1���큷�"���>.X�'�1y?=�$�Ji�5�jn��
��fc��t@C
�b��h
�S0����eq�MrK�p^�i6;�ݜ=��,�W��s�	�oZn���Iaz>7�UFs����~]��^�|�{�%&�R�����Ɓd�B��!
E�����T� ��^��q�1m���a�܆/-�+>$�db�UU|���o%U�U�Yl���3����I������Ԓ����`�m�2��F�xO�xm��o\}�\���Ƴ��ԍ�Ԉ�mIܹ]T���	4�%�H�y�'�t�9�^61[M{׬%=��ʍ�HbXGnL/&.F���z�[�ÙM`p�E���h���ѳ4��<�.H;v��1�H���pŀ�M�4�LwwO��Ĥq��2����P�������/S�L�p?d���\p��i3׀�
w�%�!A�/��f� <�N��̸G{I�%oS	e���ը��R���F��@���M�&z~~�X4`,�"�f�M��MV8�EA|V�C~����-/�_{�KH;�XppewD�F�vt֦C��,b�Z���W��WY��(kޡ���-W-" ��/.�K�uP&˔�7e����aA��T���`����� (5(��`9er5R�Ǝ�E!�L�7f�d��LU]��^^
g�6�=;7��*M����om,�B���PF>�Ľ�#��.Lw
��S�{�G���Y���q�w�-y���%�oſ��&�Իo�&��`o�������,�f�.R6j-Mع`�j�f���m�Z���VD����]�]5a����Ijn��\����kZ=o����Zwd�W��~�ۊI$��́��Nj	\��O��n+�^ȥ������-gg�u�[�7{�I����*c��^�������&����v��m������ْ��`��a����< v%���O���?s3�׼��/8�I�	,ǜ:�0{��h��&6��&zu[�Ƃ��Ġ~T�)O�9���/C�ˑхҍa&�K������0�t�A*Qm����t�[_�FE�D��Tv_���ˢ�����ol�칻]e��w�*L�m�84��9�g4��?�%���Tˋa ��LT_�"��)�Qib,*�ƭQ:��X]Mq�i$>>^����U������ǿ�xeqsm'AZ��Q�L�ƛ��M�ƆaH`���W��!e��pC��o=:m�{I��pviB�8U+�xK�'�`cmf��e��1�i�ܛ=v�"��f��x���8]ό��7y"C��Oe|_ߙ�kN�����3�/�}]������;����w3��	�	۹"�>�ۏ�`�.�7$Ѝ��ٹV�S�yӲ�����(��c��Ç/�N����.6~,z���y���N웧�K׃�Jw�÷��3�_oO��	�:8�����r�޲ԿJEEߝGT�|{Z:<8�t�����9���7�6B6����ۦ����]]ׅ	+~��z�Z��_.6_0L.{�UE��ֆO�qD�=a��+/�=���h�A�	!cW�n���h��xx�>s'P/�/��>����"-����^j���{�5^��a�^s�̯�=�p�R~pRSB�?I�H��2.����8nٞ�F��Ʀ����d�6lIU�F�_�-��k���y~~>�E@$��-��y*�x���/��w�S٬�;-�;=�>�:]{4�w�7��h9�w��I�{�?�[�~&7��1mc����|A�	��*3`dxV0n뒊��k$���ڔD{�yC�}�������"i2���;nqpp<��A��V��bL���,�F[�	����:�ё�ډgܒ��ǻJ��'q�$�h�g����Ol��SﵴjwJ�x��1����A�hT��2�<x�������`El��V<��N�w���Q����􁴹��7j�b�����:n��s��mû�<��ռ���>x���Y$#t\�+�ū��5-7{��DT�V���>�0�UH f�	�_:ڪ�ƻ��^�"$z�����QAg�W�C�/d��/��R�rBz��GCZ܂�_\9�"�2oipc��	σp���Jl�w�u\u?}�	q;��/~�������8��?!��}D�$gZS�xk����4@~��'̵XHK8tk���IѲp{�|Z�g��ҧ�-7����v�sw�ϖ��������QOr-
gn�ϯlo��[Ni�<�q�!�Z����b�6ƴ�~X��8
r2YaT�2���S̈��CY��Yt�zz��7��v�ߵt����ۥ��7�}�u2J���7�R����¢O�K�4�������-�ٔ3^�T�=�GF��n���^�#[hp�a^!%�(^�5��C���}�"cc㭡���~�%EEҪ��6f���n�J���Rd�`,;*�I@���?�\�B&����9(U2���cǿ�]�b�@�>Q�
v�� �����B3upso���8����������6ʊ�?����ZP��<���Ľ�&����:���\# y���N�T�]"+���y��D;��sW�*���2���Ƥ�Ϛψp���&�'u�-,x3A���#U�d��9��]�p�������C��9���������� �
�U=?�:�1M��������O�j����~������[�j�'�������'#qbd���J#�p��w;ZO_c����S����w�B;u�������z}��1,`�%�JI�����{ؒ��<�	j�Hμ[�5�Wn���֐��@�p~B�i�kd����6DR�#�D����j7	���&��$�頇�N�s�$h2�a�P�Ju��e3��j�T@A��7�2*/�n���@�@P��.�;�TM���D\v'4���^|ܟ�;�>�9-��BZ[/� �c?M/!."�m��~.�BV���.�
{�zϢ��sh���L�^W�����b�z���F�������������Z�*������^_���H�蛘x���K=�$P� �Պ1凌�aΈ��GuƜ��e��j[ǷP�����^C��ӣ�o�'�\_�9��ʾ��T���k���?W�Ԭ��qeju6�Gb�z������pA'���-�Jr��TW�y�����B�����a���`&��U��U��f�������1�>�
��w��$����N��`foݐDW�C�N���33+��䍳G?.G��[���G���G���ߑݤ;~4���o9���`���x�����֎�g��еT�����_��>���$������.ZQq���a� �WppN�Y�د��V{�m��:������3��㘢����UV^�x�<P�T#��x��I����]�ً�Q�R_�� �}C���������D#>s���9��V�=n��7W�xD��WξSz��T6[�I��b��=C�"5��ޫ��YÀ���<�Le���χ��&�ϴ<�ѝ/w7}��+QgCZ	-ߗ)�-\[	U6s�#����[S�D�����j�3��߿7&�8-j���*gZ�n�B���3Ȼ%�\.��3"w�=�U��	q����u+�>!SS�:!/U-������	
B}4�Yy�_�����B�=���V�U�Ɔ뛒I�h#�:0���Y��	�挋y��f����u=�j��n���M^O�����f,����\41V���F{%{8 �k���ND�>�I&T�d����s6��3%A��	
�J�l8~7m~�AÞ�����ǎӹ)�l<m~�z+G�T����s�
j�*�+�k�]�#�7\X�������.c;-O!ydQc���5Qk��w�䉍��(#F�(�V57�~6�#L	�j�~g]4��y{d�wd1��o4����zܨW�
��e�D{�e�ԋx�njF����R�W�*���	��
%��������r�S�z]��$%&`;ڗQk�J�i�1&<���(HBv��}��Uŵ�Ϲ��Ĵ/�&�����-���6*X(���F6_�j�� ��������A��ڔ�03���{�	��SM
��yxϙ��O�q��k�$������|:*�?Y	r���~�]᭡��V�Z���HP=	���N钐.��ւ�6�]1��Usy�������$!!i����H}ʗ|��>��ޚ�A��:&s��w�_Oo��9�\s �[�SGb��)Y��@���[]�����*��Z�����臫I�N"g�әz�$�m꛷��rĜّ"�m��m>w��}T�A!���Y��
X_tDɏ>�eP 2P/�X�o�_����Ȍh������L����Fo�5(zj(m�����FFV	F��5����Wg�g�0y����R�\���y:�ŋ�Â;��yoӑ��y(��!��=�zF�t �*6�0~2��k�u�F!`Ʒ=ﮖ�P�ͶShT���⼜6A��?�q�o���D�C�e�9s����.K;ǰtX��`g�.���	ք�԰�4Ro�-i�:1e��yфk\�۳�Tg�O(��zD�sW��̵\^���֋���V9�pa�0��|��ĵ�0���"]�}�����B�!�L� � <jiF���M���$��P��N%��i� Fay�I�P���M�+S�'����/�z)
#aYEZ��g�U��c�����KM�"�Ƚe�'���G���Tw�tĨ\�fv�P$��u:X��.ikW[�k�@�@���Y��o��dL�9U�i��--��kZ2���U�XC�E�,��@�Ĺ��HK�@;Z�A�IIw�ɶ�9�k�B��o$&�h>��4� ǌC(��h�?qY�{y}(q�3�r�'���Yc`8��T�$-�/�r/ȍý��t������� ������~���Q^^nZ�}坚�J���`��F����ǝ�����>���_			��ʨ��OE�E�95��U���{�^��� r�#��iO��%�_�y��9Xk�lu��p�*c���nH��b��E���W@P�7���&ꖲ�q������=����osM����sQ��C���Se�s�.QG�V�'�DF�ҹ�P�.�#{���s��`�Nצ[B��2����͔$�R+�~]_O�u��jIk1�k�O#	�����hSTr��bv�������,��S+>�$pT���v9�Q�>��l����Y�����,-"y��<��C��{�$:�Zax��#�������������տ����3��:���WJ|oI��0U�\�W�Z�t=B�44���f/{{{///^j���y!??���lx`�n(����9:Tl���;��.4�X>o!���b�G�u��b\&�#�&��4|RV�g��D�"튦��a���\�צ:���fFL#��o���ʗbM���(%<u?�9��6^ҳ���>^b;.-(b��e��7���ֹ8�.9��ׯډg��<�l>J ~f������A�K��}ode��%�*Z��q�VC�%�PJJ����˭~�?�[�K��r��j��Nm�BZ�����egg��M��Q�q(M�n����JCC#�Iu�t���dk�����z��5=?���e`^<�."  ��u��/���מ�ձ>�oȨ�\yy�O��@��@~������gf�hh�/�ۛ��]~^���2;�~w�<#Z�qs`l�oݬ�q��T;"�,&�R�]3��rT^w۷O�I������_����?��N�,ؤ�)R��yӯ��U!�\>��U�,�MS�~!�0�����p�	w��e��U���$4�+f�4�����<:SqVj�{d!5�n|����Q��<�J}^i�9�:F7a��_�:Ư R���疵�$��(��v���v5'��X�o��8���w��:k����T,0.c��C�7=�������-ib\�����
��nM���,_�al&���ߤ�*��$cj����W��P��^�Ԣϝ���ɉS�-MG.3���RX|\����Z�Ģ��^�����䴈��P����*��X���U����6O.��*�HE]�Ŕ����f�`�ČÎ�]��e�XE��v����q������׵dN�����Ɗ�=[�������:����mEA���5X(a�#H�����=#����q��еڥ���h��!@&��d��9}C��K���*a� ����́�Y���s	">uO'�9�c����?��8��jD��������R�IR����t��<93S�y�W�7�n>y�����߬eĈ:�#>������v���W��v�v0�6ݼ��i�}��b��ޞ�Q�Z3
�[���^+�-����߉��h��II�<��O���Ph׵{�(�~��b,�Pkݷ�c3�I����,�Ge0��xw��;�V�e⤀�Np@�q%
ѭղ��o|'����E�<u�j�c��R:��F�3�"��=��1�ZwC���riZ��Y��"|U���^6����+$��\����h�-8U��o�Hx���e��1��`�����.4�P���/U���VV������T��7����=ܦ��Q�JJJt➵6��N���wGI-�'�UE���,��r����zn�-#/],�Z�O��G�#̊�'���B�\���aE�9v�aY�D�}gf�q��&�l��k��c�z�d�yI�eOR�~��?��cQ�q�(@j\/O���5k$}X�����kj��<��任���
gHܯ;��9�G9XZ>�y�,����oOjN���I���9*J';lPn��=���Σ�ԙ��=�ur�Uo�,lq��H���B��۳������Z�q����榲r¢J��������G[����E��tְv�]�P�^��˃/��"�n^�WU�����F��3��su�x�e���Rur[����1Q�v7�Gg��������Y���Z}���Er�vjX��^4�����>�,+��z��㓦a��.�*t��O�w�_���ky])����0���	�	�i�B]d+��P'�����_�J4T*B5�kL����A�iqn��w|����ֆ�-��@��of@��Ȩh�̬0hk� M=��{�|
�ό����"�7�
!���v��ve�+����]����5ٚ�='�2���dqTT�X�J��yʶ66�@�<4�� �G.p���Q���}�s��w߾x�u�T�������!����N���AY3��:�z������X�M����@fuuBi��&3}}�;���U��B�N5��l���|��J�G	|u{�|H(CWp���1k�}��Y�d�H|iL/�F@��������#�еd�(e��2�_G�i\���tٶ��vFMz��-K�\v&�]��4
!�<��+A��[@���5;o���}r�+�s���߬�C`+����γ\֊���r��+�����ߞ��1��ê�ّL���HB�yK��#.z\u��r:��U�aF1��FgF'g��B+gF�Ç����$��]�M�����r9�BW�3\:���W��\VUȟ�I�Pa����}j�[�{�������"��gUL���/�)���p��Di�����k����`�?��jqt�Τt\��A�Đ�54<,q��q8�	1��#��H���L��77Kw7W-wc
/�����yTOX�;�ai��fl]4G�����7:�Lޜ-�ݯ�yh�/&J���P�(^��>�%�ܵ������sٝ��`EWVV7�=~����!����4/{��N/ǁ�<����z���E?��b�.6����j=��{���,mҳupx�n�#2_]�͛���U\�W�^=�_��}���b%f�=����e�QΕ���f9I;���!k���%q�K��hcQ\8�Ɩ!�v?	���9��$�#:���~f8p�� ����O�����,, y�]�����y
������Д�y<�|H�A�Jz?���\`�y���ܠ_�F�E�D7����t������+���<��ةT�cv�=Y�4wq�eW��_��}|�l��N�m]+ș� spd�A�̴�7T�ҙ����.�����hD���ç^'�\RCp�٢��$�8|�ai1��Y��Vu^p=Tb^��_-�X��W�)߻��86��8���n�Z3J��䋝�dB�wO?��5,��Ȇn������5��+���L*�+�x�BI`�7�ܸ��q��)<)((6��Ju��WcI�<�&g	d�+�`���3gk�O��y�����61y�)2< 9-���WTU%S�ȵ`}b��!?�**��/4���b���kX:9�I�O�,�h¡��6���n=Ͽ].�B���@���� ���\��p�= !H?z��"��m5$�Ѳ�&�HTnnM�QĹ�j��� ְ��ܐ���D��=[�+t �ߧv �<�Y����V�Dd���UU������NII�(<�o8Xl�j5cE� #�����T� b팢��A��߅�I�J����;�������p������?���t�t|CŸ)t�=���x����tr�?�5��?u"�6V05x�8�9��ۮؚ�^����R�=8�Ҭ",�o�`b��G��Bi�%���9uW%��fW4�>`����4LSU#���fy5�6�H
�f�R�H[�E�컂'����G�-��-)�' �~�M2j������'s�a����lrr����k�'�>X#y���.X+3���Ҳ�V:��S����D-WBk��J����"���]yA�Wܐ@�vpG_ ���Y��̨�-ݴ���E��F�oN���x"lj����ꓩQ[����ϟ����3f�aYr�d�	����C݌�ϗ��(�ol{зV�!k�@A�W��&�I���65_���cs����2��2ή���p�0�$��0�ok��1m���W���%�+���M#�k�j��
0����Ij)2�1�g�LOq�Rs�����,���6r,��_��N/FF����1є����s�W�]�|4e���ˉ�2�/�2v4�"*O�#9�-�M��Z���eJl~�e�����_��$L#��H%��J��,ZT�u�poz
R��bԑ _��k�;�e>_�
,�Jn�O�?5;Q5�V�f��<���d��
�2��y�@P/e�[�@e�.��TW{�w�?s��� B����L�\�Ϗ�C����
������Z����>C��/��b�	��6�,��q�ne 2j�шAWm
�}�H��M3����b�Q��QO�,�}nv�ߨ��=+�tQ%���U�Omx
�n�"N�i�?��;���[%Vk��-������N��joU��)j�E��7E͢���������~>��$y�{�9���{ι8~���\6]�֤)\��<aT��U�V?��I{2 Q�㭼p��ha��N�[XU y�9���!��+.pؾ����J�h��.��@��G�x� I��� ��I�#g+/BV��fT�G�v�?�5�K��Y��!�ߝ4.����3؝�Db��2.�
��u#�vy��V.D5x=���[�:���\�ߕ^�k��V�V[��8�/6��b�<_{,��aٯkd0�>�_|���y�M��0ƚ�T"�/��ٸ@0
�.�@��R�����W���"�^�԰�!a�'� 
�8
\�,����%2̵ߢ��Z�"ϨT|u-'��"w��?��6/I7#�&�z�w���lk�{��w��W��%��2�H�S�E�d�.^��>q[��N��2���C/z,S��C�嵿c@4.�Clmm��4����%×�G�F�H����(ڇ24myz����%	!�Q�{��N ����.����u���� �m�������-�G�<�P����Й-�11���"��|��Sa'|n�W?u/Od@T,2�md��k'�RG�r�S�]p6�^ˣ��E�+���Ǉ�p�,��eJ��s��s�N�6L����k?ǟ���tG��}�^�_YM��4����Ls�E<���-:kj���FVm�ǐ��T��@z�� �d������b>�m5G�U�@U���P��Y���!��`P_�3EP�������������"ܠ����{��1���=�M�$��c,ՕzG���@��(s�\e���3��Zq[k��	I���� 6nǨ�ן�]���l��l��|�#�� �d���<d��#���j�^��rtxFNR����f�7��x1(�@@�N�G��ֱo}���]	���>��g�eE��B5e�8=.���c;�
��A�u�l����u~=-�����=o���Dv�vN�� 6�[___gg�J�a��agW��2��J1"T�}��P��$�þpX!lL{�I��%c��C����kߣ��#�����,teW�D�9y��4.To�g�$��#d��ZT{�gA�ω�od!NS�����*����~�$���l!�q}��P����E3�aJЏ�zw���AcoV[� d�ꦁ����j~V�?�F��7x�G��}����n���ۆ��ou_� >����݇��C���x�I
�g�Z���H��:0D�wx��)���>��'̙L�{;�H��-/����5��S�'*VL�2#�JӼ� �ܔ^�^%�����{r��y������C!�H���bZ�f�R���g����X2�r?d���P�yCZ�`zl����I��]/?���Q)��Q(�S�8��z�A7�:J���_��؅*��ЧQ�5��	e=gn��LZ1����@�ys�ia}}}3׿�7�
	C{��<����Q�ڙ�?�7��I��ҌҍyQ��k�|��jؐ9��;�$4�\"_G�����,�f9ө&E��$����MT.�r���?����ݙ�q�$���N�k�sRM�XA݁Iq�R�ß80(^<�/$�%&�}ߦwq�CT��4!���+����2�1=A͡ɞ���Z7}}s�ܢ� ���!�	~�����Y!9G��e���#�c߇�af����S����Q�4c�4Ջ8�y�#��J��+T`�i>�H&=�r�~���rB[%N6����S�2O�.^^^~O��@��sxK�z�q4	�ָ�<��a33|s���\tZ|�\UU֥���R��������C��b��~����K�͢] �ܲ�(��3����j���sZ������pt�q�){e"a������o�Hq�ҽ��Ϊ�i������,,1樛���`-5)R��)ܱ�Ȃ��A�A��&/��O�p����Fq���Ƽk���ǜA��v��n��oiΚZ��&�Z�+���L� w��̟��t�r��������4{2[����=K�4gzϱ��y�j�+�{�8c�����Pg�Ҵp���s<cC~�=�	�yn�W� '�"3�M���a6�����8�8��z�i�(���<޸<�u���N̤on���3/�1����Ĕ∀B�9�V��:��Aj$]�V�O��7hح{����)�F� ;�-������5Mu/�R���J�2������Z,t�����r�I^�'�2)	�h�u�Q�� �n�< �����݁�w6gg�F@�}Yz�)��m̀�&C
����ԨtD�
��rW��z�P���lU2��l�S�����Β�o�c��r:����}��ZK5D�Fk���1���h4*��.Gv*S5*�� �d��ݎH�6���ӣ���d����R���:(����$@�j��zP�^��V�C��K��������7�������� �"rq�^�<-���i�{ݮ�av^z�>UQ�N��ir���}�����L5�"��%Ȓ݉،>'��'�EchF�NF1]�i;��� #���z>��1Ԩ� �`��\)�NV ��ݨ�3���ve����'���dT�ݓ8W%�k^{�8j��pFأOd���q̩�5��Q3�%1�%+HO����<7^�����RM��ᇕ���%{D?�hľM�'�}�M����4�3R�g��'�7�R�x-�&�b��Qbq���U�灈C��/]�鰗L?����͊DR+(�����_ 
态?Md�������F� �~:>�<fJ���X����͈�PA:�E��^�u��g��-��A��I�_��ê�_8v� �#'F�������?O�kdFl���^P(X��Z��yP��D~G��~U+��`^��f����.��6 J���y��ָ���&s����Q�uwT�yKk?�u~A '+���'`}�D�qi{��b���翎�~/W��t�|N� %S;V�LV@���ݝf�4�
�c~�`�L� �(]��ۮ�D�5�&�2#=�D�wi��vts��D,]!�qO�*1"�"�$!
t�����e�qޙ��6*�ִ%�;�y.��x�K�0�����B@���i/���1ij��k��z��G�G=ۧ��sH{^�Lu��T!T-���e���p�e�<z"3r2ҌOtwY�g�2 E��B��qD\�^���0ZÝ��(��Z,hT�vo��$�4�SxG�d�ʊ�mO�m��ԟ��ngk��*��KP�$��}��a��ۑ��I�kU���ARZ��-L�b����;I2���"GRj>��s}��ޓ�B����?�|J��Ĝ#�r�QY�SIB<�au(��*�ԩ�����iëzwe&�wɞn����=����9ivT� �e1Xb��˓����������Y󡰼���_�/�d4�Ɔl�-��X���w�#�)��?E�j`%�bK�{hKR�WG��,�iN�^��z�;�������2�r�㲳��J�Я��E��L�V���?&I�Tˡ�-ѹ�Z�p��/��{���KY
���8u��8�t+�ƥ�r7#�IP�r��Lh�����L�uv8.i��.�,6r����O�qٻo�~]'�3�����LP0^����;�&y*��M�2�L-�eH�ܵ���K�Q�p�VU}nT�==K��p�U%��PޡC�K��Μ�����ѭJ �+I��K{ޔ1ކ��◼(%��Ca1����$Y���Sn�kg{EW?ǩ�T�O�8�+�G�g���9Vv�����#dF��$�:'J������4���Sb��b�h���k*��U�0�9���4Zk-�Ţ�ABRғ,m�p�0noJ�\㊩���������A@��Y����ps�w�ژ(>Cm�Q����e�H<5�Ԯ������2q��#�Hׂ?)�Q<�%�N5�;�x���U�F,8>�G��c�w˻�3po>Es�� =d'��-B��{/�;�ẻ(0�J����C���e?M��������ru/A����Gn�������BP!�7H��Z��_3U�b�<ZZ$��=��'�5�Vy�Ul��f�ܑ/�������r6/0NS�c.�8�ѝ���5ɮ����t����G�d�-��zP��M�FA0&�k~�~S�w�~3��n����1=�zA��-����� ۜ0�߱�Sk2A��c<rCsoq<�E���6G}�f��&�1Dʖ�%-���"^�����ѓز^�����Z8@,��A��r�,�^��.�a��Xrc��t�����;I-�VWt�����b���A�8n�(��T]9�֩�i�<aox��xdee��J���A-�H&ff������Zm�_۾|���dE��X�}�:��ÿ��i�#�͇�O���q$y�V�>M�V!ů5A���k:T���k*��K��k4^�2��9F�6޾����5/@�ML��>ٙ���γb��2������<�'N��u�ƥ���v��o�dA�0xQ��L�X�{mVPG��ޓ��Mʕ0�G�'�2`��0��W(9'��BO���~�H��eJ'��%�Ɗ��A�C'2 <2�Z���+�L�o?(��=�Za���j�s�? ?!���>Rp���p��p�-��_���9	F|1*E@L�0I9V"Dn���Ҧi��ڏ���J'���Z�����HbT�(�ɏZ��j����fl�Q-�A�P�'������UK�~Գ㔑ptw׻	~�G�����p��hQ4���H���v���,�����@��2H�9Х���4ͪ�بx��d����c�yMX�K�ZV>�s�9\ߑ!��ⓑ濾{V��O�秧}���G������B��5���ӭ�2()'
�����4��l]qXw~���Sp
g+���J<~���,���®�sv�׼k�/�g���Pnyv�7������LY����a�D�ߡG������"��p����~L7�{
���=�V�+1	�y�
��/6�Hx�[��#���0@U�lю8%Jke�o%��M�QY[%�������٤�Z��;�Z�ֵ���O
>y����E���Qرk:%��`�7�"vw+�J������2%��z�+R���|��~���R	+�}ֽŔ�+�4�i�;.;��h�l��=�;� �ȰO"d�*�u�ƅ���({���Z�c9i�X"�R�GOvr��ҝF��/�/^���s��]y��T=�=ͬ��[p}��y��P�um����5V���666���-���:�R�G�V���Ĳ�Y>O�כyq�����������5�Џø�j�p��B3��0�wc�~('���}KHHP����Y\\F�D�N��;qN�4j�&�?	:ҩ�x�S����~?���*�{���Q�u�
$�`Ik&�̨�=���ȇ{�Nu��G�Z��~�`{t�M�$����
��Vs<��J��+F�XB��(�-�wB3!�!oi	�ܽѬ}��G]0:�r;=��gB��8��-)��r��'��=,@:�����X�89q_߉� ����Rd,G\f�<�E�}��[��c"[���T���ض�W;v[w���;T��~7Ƕb����]�E�#q�My0�z����w%�����,���9��ޚ���,�i�6������o. iD��)H�	>���A����6�ڦ�m���+9r��@Ρ�f��=w"����� &�}Q#�u]��i��m���o�!��M��i���Z����	����ȁta]--�6�����R���0��okR݁D��Av��k�!��dfe132�wɓwS���>�R�_+��Kx�p,�����Z_�w�)��qz[�Ǐ�A��vwG ��vV�GN܅W�}&�P�&���&&!/{2������rk�����M�8�&�;��-w�oVU��rǜ�dK�/9���UYȖ���V�K��ĮZ�pJ�d��M;4�"B���DC��@a�s�On<�ݨ-�^���=N���(����4-N<�%P(�3��4���(�����.�-[�Ҧ�ʋ�=�^o����S�4�\G{z�(����_fO�\����?\ڄS+�ဋ$�j�+-�G�!e�A��GU�(^�Q���$L��!����w�~	��d�RXW��Ì�y�3�'��f�����Zt(�����t����&&T.�1�� S`5V}Y9:h��'�Hv��}ZV(�WUk�I��~��7������Zw��v�����!{3��2~�䄨1����S��aI^�ld�BB\?�c=��cK,�[��CAQU��~Wg.����vp �u���B�x��0�o͊*WƊ��c8G�|�裚����MQ�eѐ��I3t寑�[[Z�i�ml�J�Xk����]ĳ0�l+)q���#B�r�������Bla&V�vF����g(+<�:� \( �1�!  `����)�����/��쐌��(�u�j������Y[��SP�*i���&r2J����-��������S��#ˊ��ڊ���N�&+.��T��DP�/�xK8&UM��V�����p<����I�,�V0�X���,cˈ��ME�C�2�_�eW�8TqT��"Lq��S��P��K���CO�ss�Nb+M$T[� �ϛ��>�
^U @Pu���Y��������H~6*��EV<V6�Zg0�#�������X*�\R+�Lٞ������'U+6������W�::�0*p�V�80�:4-m|��ɖUd�A�dc�]��j�ǧ�w/$qŅ넜��Å�l.��Џݜ��� a\����]���8����.pYSN��|̇1����=-������߸���vlm7"�-B�Ɏ��5��')���չ��K+�T�9%���^�92���)@h�+�WI�i��P�>�&&&��QV1G��m^ 1�o9���`��ys���z�m�-�v@�M�ɓ�;�hn�ME
���W�u���G
֧�z28Sk��	�}�����M����S�K�7XG'�'4oj���_rۄ=���Zl��]c���)�[ܑϡބh*S��M�v�O ����w�D��@]|�����5���F�\�;lV�����4�.�����,���5����.j�xn��|Y3!�\���Qj94d 6�l��"�}�?�
���Q�� .�/�s�&�i��0�:���e�����[��>�z��.7�s17"gקL�[p��#��"���*Oy{�ÄV5�5�ꟻS 8[������S�&��z�~�ԅ����}U�'2FAa*9.���	>ۇo��1�S�(��QQ� �JG�E�wpF��b��������G�E�[`���+�e ��/��Ȩ��o>=��A��va������պ�J`nv�1���tg�C��zF��=[�?�'`�9�8|�߮����i��:4�;I�l��ϟ��Y�-�n��[&�D�c�{o��¼�6�6Hkm6��F�|؊�R���B�Rk��a[g�&p����ht�j�>4iw�s�W�@�%�fLge�Ӣ��fW�I�f��c
�����a��{�����x�wi��o�bӂL�s����i71�oS����|�w�г�-���_cK���?����ہٝ1lr�xBR<X,#1\��R�h���S@�ɠ�@)wضtp�'y.A��f�%;��;D�a@��)�j{�j���G7�'��η�@�� J� ��A>��r�|�DU��Ô�0³�Z
�P8r�EA�If�iڄ#���6�tƬ���%~/)�Y`���p��'����/����|�Y�7}i��&��c� �]R��=:;e���4H��Ŷz�w�w!?08�̶# ��� ����N>�v�E����쭭׮ϗ>~�x�&���+b��������g��Ng�,+�Ĥ���7J� �5���e��GU	h��,�ҫBde���*���	A��� �=��_�����n��.n>�n5A�_�VK$nnl|�|�r\�\��m�ΣPP���R������;���>�`�(a�CNL?�9�Մy$'g��]s&s���灆�� w5J�F�w�,k$�
�9���b��@8_$ڭ2�DL���l��X�������߷�%��@-�Jΐ8��\(#m�m"�̐�̠��<���m�4�ukUUX�}hCK�KoJ�L���ܘ�=;� ��1cө���)�y��4`��(7M;%���uҠ�L��Խ�\���>I��ř/��1�I�e���+PԷ�`�z��i���>
rFtxh��N�Z��FXs��)�����M���:����SA����C	�jO��c���� (��'7�O�
qѺ��&�8=����8��������,hj��R����ܤ�ݒ��s�$���Ѽ����� �u:�z���<R��2F�-6_�����q��NԴ�?;;+t�\��V�����Q��9/]]�a�*�W�4wZ5���T��� ����S�*�:�6�knFϬ"C��&f�����dg��Ⱦ�@�Jf��z��m�7��y��	U}E�����)�>%��/����p��g6��Qz��d����Eb�(5�������׫���S 4u�+�t�A'��j����)�vs���d�'A���S vFW�i�1a��d�>����4����W#}�u@�c�Ǭ/=P��T��5j7ʅ�`��>
$):�g=Mb5�b�
)Ĕ�F�c{��_��;00 ,^a�S��Sb@'L�m9>((a�+&�	?3 ��r���蝳�x������K�N��<p���}e��e�֕9R)�s-D	���P�����vvE����a���F�����ּ�"�ʹ�]���x�i"�b[�^?�.�5Q�G����%J3�b�6jZH\3qBc�ӷ(0��������s!��� @J�?��-�ܹ=>����J�����C�~���ݗ��0�y�n�X ��l��\a�{��톳/6��1�K�����_@��S�����Ҍ]���Cݣ�;��SS��%��~�~~���h�����'n����� _���ѬL��W���'�#�� �.��n�ꖂ�(�n'�G���אӛ�p� ��j�.w����T	t�PAR#��9�
$7��tJ5�e)}�ID�k*׈�w������V�f��
q��q&MGv�������e�BT-S��O�Uvw��;.��K2�҈�R�ֻf���I��N�yR���YD˩+�����q�=�F�4���\�	2��
Fa{s -x3-�P(x��ɐFU��Y^mY�=8~1D��]�>VC��5f��P`z�I*����./����EEP�5������m��u��o������z�欎���E�4 'Ĵyxx �1��7M�S;�5x�n�� �eeet�MU�����yE�wG�aď��=����ٜۦ�ڈ9�Ж5��`>G�*��+9�^�1o����[��i���)!`�#��'&\+�i|S�C1}����� �ž�N��a�0���ӵ$�V����7e�9@�ו��������0b��ʥ���<��^܄�ɍ�T���G�����b�~Ծ�ƒ!��@"��ܓ'�Yn�6��c��o�Dg�`}�}���-�1*�!?���VX��`f�d�Aap��挄�y!������S�2=-�f���^����bo�ؽ�|�L��BsY�J#��1Ns����Ա��Y��Ӎ���UC]�a.�L�������4JkQ���8��8oSEq����%̛M��/��k�i�*�N8����>�~%tr����x3*� �1�o�h4`F���d�p�*����X?�]�T6���UT�I��n���wS-���:>}�n!�}��?��l-�������%ICKO��0�,���-fP��¨�oZJ�Q8)��'��iii�7q�<kċ�xa�`U���|�o��c�ԛ���?�Xz�H��Ih��u�Nm��Ƌ�L>���X���fbc��v{�u�"��x�r���T���
��@��w4����������N��ٹ�=��>f�ɯ�P*���^��{��7��h���k 
U4�cxx���&�yrz���us>��Ё[��)�ze�M�:�����p��܉���{���7�����5h�3�V �҅ϱE7��̿���#�,����z��=t��g�e��p�����G��N�=�C�-�`$�ں�k�+���!˾��"5�%�`Ѓ�ޔT���W�eA�1|O_���;W���ɮ��_y�X�$5%�0�G|�<�!�̟_m�F�=Xa��+^P����Fl�=s(8�l��ކ�v�2��O�?I���Дx�o/T�0���� q_�[Bq�������b%}��~ar�q� �B��b���}���{Bd����-��H�b(����2>G0�0~��z��V{v#�������bf$�{�8	CCC"d�H{D�O\:���]`�
7�o�[ke�~|�B�;	���a�M�G��1s�֫�"��g:�����e��U��0��߿_�S1p;;�	Նg��0������/Z�O��v2X��a��{�]]������y!Xʀhb$���d��R�`D������4@�+����*��M���jO(���O���&i6�)�����c���a��L	���Rus%_N�`���������.K�cx:!U-�H�E���AEr��y�R+���@�k�ق��<�vvv��}�oʬ|Q���p�@:�(��_^����c�B��2���VsͨU��CF��flY*�c���D�5���4s7�1�y2m�,���
�Ћ�����͐H���o(ݯI�q|C�dA���'���������"Ku����Z��t.9�|)3@j#���M3g쬱B��|�E��ǈD�W����\��j�")n���ϸP�l���� ����~�T��t�6��{�<�HK��]�Lv�@���l/� {�p������[�����������t�c#;���P� �+�}��9���!�_nQa��}y���H&ak+�m"UW�8�]88Qa ��某/Jd1!ˡ�Ui~�R��[�%��L�pb��|��
s��Z�f�;ꦞ��BGW�	93E$EF꾗��2eK��7K#�c))8r�@b�:u*��:Q��C�K݉�{r>{�����T]�F�-�������߿��Uݠ�T�ૹ�rsl�/j]Ŝ)��f�~���O��K�b8zV�|V��H��Sk^��I0+�ȫ�ߝ����@�`�����[!��%�}E��,}wI�X}�Ӯ�+k52&��SJ(����":��;�H������r\kV'~#y��觹ܐ��~����s(Rl����a&{���xsx�/��3ۂl���ִ�U��)�[a̩���*�T��F��\�0:��3�I�nd��V���0����A��I]��qk���ma*�]��Yx���bѸ��=��A�������(J	�6*E�}��5�E#0��:^�ݳ�>t����S(��_�z�M�G���=�:|!D�D�	�O����T�"��\\\mWCn��ɷ�١� (����ʌP�VM�����T|�f���-}�
qzu��K�v!�4�P�֊����A�}��N�������օ�%EEǜ����	�Hw�=���4L'�����Em
�����2�+��%�����Z�t7 r�F�loo��a;� ��p����w����h�A�US�US�Ez��͋�#�D����H�U@+�����bwY$~�y��e�4������������")|s|B�I�Y���iɹ�7���K� �G'0b5M}OΕ.֪@P�l�օǃ�.;�H|�g�s�t�r!ݬ(&�.��ʔ[C�vFb�G����D��/q����$ܛ�_?��g�N�� �K(Z߸U˧$���AuSt<��l�r�cAVĺj1�#`|�3A:��v�TTz��Q[2��b�c�P�����ԡ��_����/W�9"`�O����ַ��� Q����3i�ۛ�gϞup�Z?Z9d��-���
���W�/D�,=��~u����7贽�������{rC6�����=�����`�06l*�9e�����k׺�>�([�q����ܬ,`��h�G���r�u��4�0v	@� "��ӧ�N�8������A�}R��}ꇀ욑��h��-j���#���kCY���4ۖ���΁_qBĮI$���� ��Ç W���PغR�1[���[����vvv{�]9��e�L.��^�����[ݡ��C�J�ӳ�%F���U�N�)����neq�2��#�\�9�1��8����Y0�%t�P�J����t B6u����a����mH��Q���%�	���cZ��2�w�����\J ?~�$�n����� yy�&&-�]^��ޮjڣ�Q��l+Њ
�w�5�j�-�xߥ��$�C��U�"�+>��u~��WޫL���*D��WFV�v��w&C�=�G?��F�Ul/�ؾi0���o�1�V{7���(1òS��v�s��T�[��kr�EO�Pڟ
 �HUL�Qz��(�1������&�1�Y���=�1��Ьe%;�X�CIr���G���vw�>M�c7�2�Eփ�@3�/�)R����Ӫ�X>A�NL{�%l1����>��O\V�7޸�<	��i�Ý�0��>.�LS�'+&/;,}�%u�᮲���C�ʻ�S33�� L� �b���hKK�oC�)M䛻��َG�^3E|�U��P��Wϣ��6=e���O�\ 2:�2����u�/����v�}4���Y}֧`�O��-8��1�M�N+.�Pv󻽇/�z	p^�� N�cR�I�d���i�@�Y�=6��D�����!�5�3�&L�g���7��ʀx}pS:�Eb�"�]̑ �9w�};O��`Q��*Y�h��%!��AaM�ǙG��D��0'�-7E�����4�U������L8�%$��4�eR[���c�x���P�@�xՀ!��l ���3�L1JӺx2Vo(���@��/VNR�y���_a+� ��:%��zX1���*fr:���������>�-���OfK����6��>?<���il��Z���G	�0H��/no���C��Z�ݞu�C(��8�2ΙW�[��O�0�u��)"��ɽL
A��'o���'��ald�){�dĵ=L�N;F��ޱ�S�^������j�Y�>��re�{�N鱺Ky>_O��w3�m�z�0gX0^����:����]�W8_Ë��|�8׸5*-A�g�0%&)[~����P��xv�����e���~C����e���_e�8l�$�qaI�e�ظ�C��ZI�Ng�͘���[YZEG~�)2$2:r��2�2�2��O]��;��}(�lA����l1�M2� �ħ�U��X��U�G�/��>k�f�:������5s1j�_���];��N��Ad���U�PR�o��@^M%�jٮ�*�w���:QH�S�71�C�¨�h���*��ڪ��{ׇ{u�-���i*ޣU�;�h��1��)&_c�w�*o����x5����]%����`��6��0�A�]|1��Ns�3'��	��,�Nf�*55����y���SғgN{^Rߨi��2�?W�(}�a�NF�I�|(��o��A����X޸<��w��[rS{�R#'Uo���e��6�[�篷K+n�{]���'7Wk�k���V|�a���7�S���M�WG>2�IG�����..G�Ǘ���L��-Ѿ�ỿ.�<��p *���1�������atro�MMh�*��Ĭz��
3�Q�+Ŵ����Մ}&��'�䋞�����?��)���c-߇$DG~&��D�d�i��[��˨JI�̜1	?��b뗰{��X�~�h���M,@*�U~��QOFff�]q ��cV���Jv�H������~a�^y��(o����#˵��,��N�1Žg�_��+tR���y?��!���B��~,r��%
	}��o�Ը�Uh�dAWgu����V��/ݛC�Ց��ɠ�� '��_s��`��%�������x��Ғ1xR�����/�ݕ%|`L\@�am���w���}i�xN���/c[%�@U�����l��4��Lr&5����=���!s�7�t?@�7�Aa��U�f2ͦI�d�Zo&����h;.��RVQ��!�@�qҀL	4�����ϻҦ��cw�)<6���-��0�0�.*P����ޝ!�� #k�G�a���v������f����3>Q����Y�Pzɡ��#*ݬ5�`��{=����2�����WT/I�'�5�4���uj_~�Ո�P��}&qܿR�,$�.�1w�.@���Η�.���w;�%	;���қ�>.7�N�X���I$���hl���HO��i�)�<�	�.�tp@�I�$��)JlF�����9n�V8���7}��hl��X�3#�7����
1�����n�%ʈʬ��H^���ٺ`�|�,b���<>T���3�I�N�0��%iy���9���'uuu�%��4�/�B�Y��s�
G�\�P�Ռ���U=����v���*4��3��	>��R�D��$��I�D��B����GK��b��驤�����<��~�744M�g�b����#�.��\�^|����{;�+������r+��&�aҰ���B6��-���$�i�P�V�LU��F���ۘz�7e��t�Xq{Y���*+-N_q��ˇ*�L�rkT	(��A����hШfee��8��&!4 J��4�h8��Nnii{��,m���3|{����Z�O���l����`�ܪ������tu�?�)�l��,I\��]��B\��͢|��X�i��Kf]tm��3���$�	B�Ssy��|��ncj�����w��w�c�(��z��1�����-X1���~�a��
�s�B����x�3� ]�̟�����r';��b���V_*�/���ǆ�w�:��ɢ��}�l���"[m���Q�ǫ�=���B?4���G'����}���*���h�8��������`�A�j���BT�������b�6�;K��|B�&3�क़?��v��:$�����'?XUVRr�� ]���_Ս�a=88�Ga�%�8�U/���:��٨p�1��+�O�3�_�9Pe;~"8���"���֬����  Ӑ�#/���6��b�1�����P��0#6����O�_7�T:�=�s�a��L��}J��l���ҧi�V���4�q�]c��K�pT���ᰉ&� K���^�;vh�/�K�9ْx�ͨ�$22�6����F�~R���yW;K��F! ^iu_~�%im�$V�&U��R��9�JOʁ�MJ��@��ܱ^���$�A?8Τ�m�O�$��׍�,���Te����j�U�Z���-��){'F���4D�|����
��ɓ��~n)O"�ɘ�<��:��!Ԗx0����c�W}�D�o��eldjJ1]�O[j���+sDL2���d� RU���[�L��b��U8[�X3��W��e�}���{CwU�)7h2<*���ӳA`�{�ԵB�y�`��_�Eֿ��k2�?R�"���ԭ�1��A@�;!�k C �ǚ��=�yP�Q�_�D�H����Ɖ���ɱ�z��9;��ػVRR[[;<2�"��G����P֓H�Y;�+3������72�z!�!��,"w�_כZ�z%�i+������������`\)�;Kw�j9�k���ou����Cn)��	�������A2��#Q�H�Z4�H��|��A7����t�jͼ�Y�'�ʌ������m�����;�/Ĉ;��k������TG�aXh��Hl�5�z���i�b��jZ��0����N��/'��~[�;'�"���%���oy9j��������u������xj���Æ: 0����Zˁ
�[���=���j�U�|wr ��,)JcV�?�ƴ�n�T	������-�O�)5��	:.�:+��M������^��#��mR��Ʋ�#����~�=�ȧ�D��*[�H��O
���x@�Ĭ����C��&K���I����9Oj,�j�@z3m���+�j�%�q'�7i�uO�����_�b9Rx��_Ə��A=���h�+������[o�� ��v^R^>xポ��f�bg��
v�kD+�ֆR]Й1`�o���J�o��;h���ۇ)z�֚��Y�d�v�VV�覞���z*��qX��Q�V�Sd�������8)YR�~c�w�8�;Jf*��Bt��ྲྀ*��S8<��n�̨�k΃7c�H�ŋB�������d��/'4f�Q]B�4@RV�U�����{��d����T�ٌBM�~��c���&����&��I[���,��������2�%����^��7�)��\(8ٝ�`�$�+��?|�+��������[��ө�b	�-�222��*�^����ː�+�\���O���46����R9�U��iF��bqrt����-�������&}�Ò�u���bq��$�w�9Z�;( F����#'bکg���~ 6ɯ���~)-��M_�V�t�R�(�@p(7^\Jpwwww��ݡH���%Xq��(�X�/<���ɏ\��g�Z;3�j�D���^�UVU���xy{K��nll �A�������Ի�~�C]_K�#%[��J  ֗��B�q(fk܊�#�N�p?��b�Hc�3���H���MfH�j��0�m�@_���`V"2��;��(;F�m-Vov���v��ravD���i�3V�F"?ۻ�~H�/\�B��ć��/-S*��ﭫ���ԧ9�*L�p��l�quf:j�ײ;�Lƣ)���R����-6��g�	s0A�J	he��XE��l낎'��C�oW���̮����E�z�p�O��I��$�I����\���nt3�O2;����]�A(S�kA ��3���<�叡��zۜY���	�����E���A7���������4*���e#jM.h'�e�2��b�������s���҂���Tߨ@���7N���?�|����]7:J��E,��^?�$���B[yDz������g���!�w��������!꣢z�鿉F	�zJ�A7{�`�!D�.�p����".
�-u���>�3@Bڨ�͒������͞��4躼�=y}}m���#�^�� ��Y�y}���23�x��R��S�W�[���fi��(��ڡ�.-4$�	I�͆�G[ ��j%���J|Ći�G3j�)M�
���v������̵r������y6�0��ߨ^�]�)�J��K�b#p��p@���F��zD�~�ԂL����ur��9��_l$�jJ嗛��O�5�k�呉�Q6"���v�v_	�d�I��������ƭ��),  fk�|�H��/�W���j���^<\N;;:n���ɕ��ī ͓"�6����/e�G��3�Jr�]C��c���mC5ZY��2۲&[Uǝ��ƫ��k��ل�D�e�� �'Fo?��� j�V􎪪�~x�cSS�;��Լ�^�;+�Lv���/�ب.��A���0��6����o(�U������R�q��S���dZ<�+y���1�
������W���ݝ/����}yy��%����P�Xb
��uY3�SV�	dp���~l�d��1[�Ǆ9\��(�*�xI�( �JM�31��$8G"p+��L���r��@�9c31�����%7�+�g��#�j�Z� ǲTG%k�+��b-����b�v�iEI���EƱcX�љ��&A�!�Y�ȴA��5SG£e>�%4H��Q�n@i���D��jW��b��(��$�y:�����M�Y ����Ugm=FS��,c^;�U8���x��"]ܿ�Q��vT_��u\�Xs^������^��!4y��d���(�n(W���8�c�7MJգ!�M6��6�]o�ZT�Ǩ�JR�Ou��7�����J�*EI��11�*��oB��K�F�<_B<�h�L�
��,">B0�b�8�ʊ�\�,�E�x{�y��1��W��y�������WMS�,���(===	8�{��毴���B컿}�ťz�ߌ|�V�3ꎡ�1 � PV��k1�y{nu1w5�.�i��]n���X67& ���ɫ�j\N��#֐�\-d�X��%o�9�7�6��?��pc�7[T�c}-��7������k��
��-�G�c�Q�FPc[q������aY k�T,�����`�Nk�bV�7����@�V	�܊�E��4�<:�#��Ȣ\�B��(o��F��n�i�[P��8g9z�`�m�g5��3�u3�lK�7[��4e���3�L�,�}x�4@��I\��P��03!UU�;�HtІ�qX0�6z���tߨ���HX�zd�DS�Ƙ������A���6����|o]r��2�yG����	�yC�{���H__dd���[���E�ʈ���F��� ��w�c%��Bʯ��sy��p���G�~X>Җ�/S>�������-�Jnn�P�߄[�N�����!�ܦ�N��4�W�Ƨ1<����a����5����3��:�TͪJ�8����|ߖ×,A�h�����[��=��\�4(q��*!��~ Z����,�8 M�U�`qVwI����]5i8����84��uB�:*�H�۸��.W�Y#^^L�`ۏ?n��Պ���J�!��|�(�f��%M������	ú����F���.4���*sR��A<7R]2**�~l�[�I:��S�&�&Q�pYc�j�W��d�&��������� ;T�O�
�3X����M�4�$�l��	$�Z�Z׮|@�+k[���a���f�>��=����|P�:b�m]ه������������'�8�Z�E�-�Ӑ_�8��.�����q|s�qa��l
-"T�[2AlVۀ�#C1�e�zTKKK���P�(�#�e.�XV1A����kkk�B�0�p_�7�5a������Qb=11ѿ{����p�0���N�n4L�~�\*䦧��[q3�e��$���Fnɞ&�oa��u��I��c	n^�]N�����w��9׆��#*�4f�M�o��t�v��f��Zmr�UĖ*�l��(M_>��s,,#s�0՛^Eiћokm�k�Kx�}��C��#���"?��w�荋��̂柤vCH&Ԙ��l�t�#�w��w����s)4�b�ݗ�c�tf�<"	�;� (�b�$��t��j�$��'�(K;)Uks�|����|z���%�_�S���윹P�B�Fi�?qh\f���K�����g�cT��e�AU)0�C���2`.��'��1����.�tI�����@�S~L'%�Fn��W�XE~�����*����>�a�cȦ�`������!y�.@�m���O��gUU�����1>j�O��/kz�~�%�M����٧�j�k���"�z�d��g*�gb�EG��:��n���:B+�N��ݏ�7�Z=!��'���8vK�6Lt�����p7n0m�ѥ����n�����㧒�C��c�	�P�<��j,��M��ȭ��w���tt�4$�?{�6��;GF�;�KB�zc�r���Q֬���2�$��顾�8�.L)�q-%
�Q��d0²{^��[G�uKrL���ps����Ӝ���u2�M���-���gK'���bL�3����F���{��C����M�骿����e�ym�]l�3�xa��OK��pL���J�z=��p�E6͠p}
�"NP����� ǭ�(�L�1Ѱژ�B���]�?S�Wt�Z(S%� ���~}���(i����Q�����x{��(�ȼ؛-�͋��/'�z�-�:Ip"wΗ�aǺ{-�KQ2L�cf}N�)���3퉧:�=�(T�MA}n�H9� �ry�%`���^���Y�OGD�����_�zp�������] ͪR����S����T�E��|��Hf��*��͞�Ƌ�Yk��B�g�y�}���z��f6UF��M�C�!?4kPyh�ƴ�X &[��= '6�c�Zi����X@�2�\�����:����z̢���9`y���z9�J;�(���JdV*���!7',��>��yj�	���������:���@KYb�Gg����=�|�N�p�k�K�&�[�$sV�>����е��@oD̿O#��� �~RFC58#�c���R2%BiPy����A��`����(�$��.>�H'NY8�jc�(�{^���mmn>~K�4~�)W��NH��楞|�G������/vEd�R��	.�#;B�G�S����$J�r�e�����c���/�wF�QQTf[_�Q�iφ{�D��!úgPӉ'�P2tݐ ܽv�_�Z�g�kfH=}i]���<U[W�:�E�=�c����2�m|���w��c��h���y���ʿ������Hi��o?+i��v!Iddd���o�-� � �o:c��U_��GP��#LF�b�h>�����nbX-@0�$i��c2�����V&)qk%�r����Z�nC�b���B�d'FBC��S�MC����!��e������=��n�o����>*��ܻd^Xi-S��g�:[��uigt��|�]�a��j��ǆ/���	�zT�q�)������}�ߎ�D0�X`Um%ؔ���>l�}�n��t�q/�X�K�O;y������'�K����n�]B�͉��S7��	)%��]��]E�u�	�S�2>��f���B����Q���>4&����i�&x�V\/���I'�R����V�xf����]gTs���<��Xh��M,�z#�]��^���*$eQ�i�W�΂'�#����V�V�^@҉�dT��n����?M�������9�]�o�On�~
�q����k��ך2��f�TJ��/��n��.7P����s�bG����N�r�����m5���ߩ�]1�����R�׫����$�3�;328t.d�˅����%h��2�����a�`:����qP����Ĉ� �l�/�4JJd�V]W�m�� �����jr��7")l�����s���ǖ��MЄH/]�iyc"y;�:ٔ>�R��):I�7H�4����m��-���/��,�=�>i��͋���umUI�L�R�A�>��r��i��z�M�-��`��m� ���G2Zș^�'x��vg�['`vu�����O��3/l��V��ȷ_U�s[�(�6%���&8�R�-,,�K��6cL���H�˕��ʖk�R%��χ�v64����	)���uuu�߼��=���������ݞ���q�������T�)C���w&��%Y� V�H��f�w�7 �Í��,Ä���bD�g�t�A�<�8�����ONmG��#MUWD}��u}v�������i��a�W��(_ax��[Kv����t��������N��0O"�U�3Zm).pđ��$��F�iP�.]S ���x�=;iL���t�$� �wz�ة.�@��ܠ-�F�b������g`jN���ʍb�KO����O7]�l��r�W� ����(Ec1ɞ4��^�M�c�J+F�$T�Q�rIEҮ�$Vhq��J�J���f\�&�e������ ��/0��'N�/�����z�i��t|�:���镧b�8z����s̒��x�+��<3J�TY©�*٥p]�e�^۟�p�>>������x��rt�o0��&�J2��(U�[H+[����9} Dqs�8l*m�2d-k��Ĭ��|i�2����K�34MSf�ٶ�'�ɢwSy�;��Ez����3�K�.q���|��R��������C7�ˇ]����+]�<�i�ٝp@r��qb.�6�\=e�M�If�&΂��(梊���,�k}<ͅ���]�l�_�Y�8 <��C���W�IY	q[����(U먶�A��.�CΒ���\ق��Y��%��tL��^L:�����}��9K�W�p�l�JKL�J^��`���Kɱ ~TbI���諿��M9T��Rݴ�ǐ�2�q����a�̄�k��k�����Х1v�z�����- M�'�X?�7.�c�mʹw���ǝo�ؿ���j����HL��i��WK����5�H�
��
Zw�w����l��x�ѣ@�h������P[���e�&�RQ M`����3���q&����c�{�iZ$��>������.j���
w�bg�ѡ���G�ߗ���*L�W1w�x��4	/�VVH^��ݟ���>��P�(^lhkj.�����uG�Y�,/R#)ן��{�����T�4�ijd��6�W�'���۸�@ B�~����:#F�'~ڴ5��o(��D�5�)^O��#/M�-)ؔq2�:'���LPa~�w<���J��*'�A.riX*��@w�C��iNƱd;�!�щ��$�yp�L�[W'*b�Qg��t��v�j6L�o;$�k�Z�W�.�����Й��K���M�tVp]o�P�Kɜ�K��V�h�G\���QQ[���"�K�]C��_'��ْ�Q�ջTp�D�6lav��p�#���V�)���xCp�/��
��p7�s�Eo��}y
��r�rx�sO�?ȧ��t�hC�ݪ[�2d��-@�	"Kc�;;����NlDU�Y�:�2��!qq�e��$�5Z���1�nI�5S��ޑ@��߻X�p:���ɕ_"��Q{��N��סd�N�h��-���p1��b�#�9�!�[�մ)�g��ǭE�t�댺s�.�ߵ��|md���&?U������|5��\��U�se9��j�i����������|
��5�q#��F�X�Q�"�*��Xv�a7j��$���W����IŘ�Տ�� �Ü����V����7p̎��������cę��+���:�@��&�?�)&���M�����i�5����M̢Q��m�4��L	�@B})��J++_���ÒϜ�l#l!��I�с��NJ��Ö4�,��͇�����3����-
�j�ι�����_u���+2�]=��i�%��}�rZ��@[y�)�ƙ�t�(����#zۏ˾�!�6!d��Uf�2��F��B���E�X\;��f�����yj�Z<�|�x9߅/|�M/����y
"p�y<�-��|)E������	�7k�a!r%��Z���:���N4n�� dR������u.��0�*�s+fX>���;:�M��ԍ@��Xr%���H�r��8~3;ꎴ���Ⱥ���|7�����ĠO��n�m�5s��[a�ٹ�kZB�,����ߺ����.������SR�c�dP�.�z���U�hjz��FӘ䋸=�r~��<d�({��X���+-����P�JA�=O�ݷ��l�_Qx�L|ַ��6������[�_�����-� �2������`�>�l4i�G�-��,�j�ݨ�A����C�w���j��Yh�$�����I�7Ō�j��ͥ��|'���_l?@��R�w������pE �d-�#�r�QÒߥВ`��t�<��3Y���Uޛ�(i��G\�N˙�~����W�M�f�#��k.8�DI�&��e�JFhG�K��Cᐫ�	u���c��֞����ѐ'$4��%���W�{y���{�.�)zk������?w�ъ�R3u]�d�2�%�5"Z���Q]����ΰYCCCQbGO��/������أ_g���,j��5�E]__���1����e>F����`*�X<���r��ndS�����r��j�$S{n�{�UU�kbA����&^���,
3�oo��5�Ϊ.��MY�Z��iG\VV�E��!y�f�r�{�bx����B�xom�|8]�HF�o�k���L��'�� ���k,,��M	�Ui�*I��������̹#�&*��F�R�����@��9R�1���}����އ�����B@���I�"��G���/�zo�*���ʲ�2ՠ~�M�T/��d�K߁�>0�KG�v��:m)�t!O�u9��_N���`��٠�����������n��J�#��ߞ�Ҫg_�2�d^�ss�9��{���4M転��Li�FC�i5IM͟=����}4%!��f��R���.�˲�~�xǮK	�y����OG�W��_մhɚ�L���V����Qu�B�W��jZ���D+E���T���/.L��K���x�.G'�B;v~~�P�m:,�i/A����w�-�z�7����]_S�_@�@���=N��!�$^�|V=�(Ǥ��S�������Ӫw&�@��W����he���q��J������;?�x���.�Y�����J���89�u�eQ�ne'$��-�!��Ņ�/�=(Ê�[��<�v@+';1��������c�8 �_j�`��`T+�G�
RŢ\�M��H^=�E*���*}܅����Ԃ.���B!9+ƽ&g[6�ް��r��f��}�s� �'��::������Ђ���[>��2��EdT�X�8���UU�L b]�6��w�HǛ/����c���l����)//_.<�`�M��-؏.^:�~�w���[H2�6/��4�]���iZq���yz��;Zq��(]�vG�����T���̠��ϵ�DJJr�X����(Λ�����/ ��ex��!I�sڵ�u��Ϸk�O����-o��k�����F��4~�v�T����HfX�����Z5���p܇q��Ŗ٢�!����ɍ��16y���="�����555[��Z{B5��p��44�̨?��ښt�45~$�>���a�������y��V"��'w��T��6uw}�d�{
��<��!ߛ8�`$+s��N&���'7�V		I��=c(�ds�pA��q2f��9�c ^�ɠ���������`� �7(��+�N����x.�xSe���>j!rqw}?��*��U�����o�zjr�j5�	it�]�1�k��s�;yĻ��2��{)�<�9`�S�M�:V�UU9�Vਸ਼͠�����#&���������Ѭ�GtР^��<�bV��%'�2B@�۠�*fD����1�|u/�/ad��0���!{�+��){�!S��m4ݦ�0������1�#vKF��Y~��]���f@��H!B������S��Jq��a���$ak�%$&6�&(��vΡ��f�q�j=Yk���	j��ۿ�L�K��aϝ<�E�_�_��ܒ�ؑ�UU8����ï�K��P ����ҽԇiτ=d/22R��R��#,��[q�~r��\|l,���di�g��!��Lp+�r�WlCM=3���g=�#  ��e���p?I�d��h��I\$#s�$��7��������Â.�Z҈Nd����?$)�v`�* �q�dP+cl��,]�e>����<�}6U�6Ə
�o���_G���bBIb�ʴ�|]Wc�f�{HOVJ�V�(S�x �0'��S���/_goto��)yr9���:����P|td��O�2�v)�ʑ���?���̞�����b�y�S���h 1܎^v��o�d�òeu�D�ye��T�x>�����-��@��f��R%��5�khMVc#j"�y����	�������������w�`4tv@�Y��[���xi�oj����g�$��0qd���,���ᢿ�߂3[���`Y[.���4ۜ��=7��_dîye�7=�G{nw����hY���G.�[�GK�����Ӳ����U*G Г�~U�\
jf�~��;p�ۿ�eB����fؕ�;��!zn���9p�S�>���!ގ�Q�8~�GY1��v)b�E`����@��9�v���K�9H�F���Yl�	~����T����H5_ sI:ͼK�am�ȟPڊ�g�YC�̥Fq�'2��1L�ѫ3�2����|���BR�$��a����Q�"Uި���Wu�Zk��`�:I3�E���������)Sv��Lld�-��퍩���D狋�onD���f�p?4�{��ĳ	܎�Pv?��w�/u�PCW�J�Բ��~yu""�5i|��뙟��Kz�]������h.W�}�WvX���sU3���vc��uoo�(�����:����1��Y6����QFT�����X�aj�z����
g?x�x����h��<[����ٸ���ۻm���x��ϟ<0	U���bP��.��?ډ1���(++u¶�����1�;�J�ʺ7��55z,�[3��R� x}�ufU0�0���L�*�_�M��ɵ�CY1��)��V�ɠ�����R�	�㱞���ˉq�T�'r�O�f�&ƭr��@���� rFgM[�����ވDC�d�"I*r��-��W��1F��/ MX|���b'�Y�髞 X l�Z�B^������*E	���+����POytT��Ks�+2���A\�s���sZ�a�F���մ�xvX>E�]eL�Î�?���a,6����^�giW.y'uW3sGKr�����X�|����T�
T��c�c!��-��H}���~p���m���tB�-��=�?�|=��/�7��N��r�;��%aa����h�����`2L%���R�dQ3����̨��3��^,Y�/��&L�����3��l���5�K���7?�<���$�>�{OGt����\�ڙ�P
�U��p?��O^Z2[a���B;��3���蘏Xyy���wï��,�dߗ��@������e�����0>���o�л���OMO#vN�Za���'��0��a	n}��O\�!�jp�i�����峼�J
�'`n�H���Q脥mܫ�W1"}��������J��#�����\1� L\A���Y*x���f!�"�iis	��g����5F�vU7�]�9��1��v��.@�2�[X�qydNγ��5]���F.���Ll���ԑ3I���E��68�#�0(�]���4�5x['���y7�S���L�RPJ�<f�3�ԁpg�}.i�w�2l_�_,�똴�v���[O��k��ׅ"�K�A���G������o��C�d��I�S<53Ψh��xLАP��99�u9�|E�۬�ʬ���R��x����w��A��ʢa�i��(F8D�1��t���j�$�'!ї���I�j,}���`�[DPG��G���f ��
����[8Ͳ���i�C�>�H�A���^��=.�)�)�����(��w���f���� 񂤘� ""?xç����bM���� Գ�C5��r�_�V?N{��?�p1����>.�H�t�S�/]OtLE��vG��9z�)QD=i�[��4�tő��h�c�$I��' �u�ÌƠן�����!�ʩzԞ���@4/J��߆�ߍ�+]6yh}
�A�����r�����<��g��-�K���߼�	~���ְ�����\�/ᣣ>�?ە\�g�w���5;έ����:R��!����#������I��Xe|�z�)��J|>`�����Q[m��I�����v���S�9���l���#�VGR8���ĝ�����kZ�������Rp+��_;R��m\�Y�skj�S�;�e}�R��%�T5��DǓĻ� �*��kc>�2���%<��8�iz���d��'��L>��AB�8��m��xS��;�e�Bv��a	��3��2�3�B�^Ű��Je��yF���|�@��ns!ƌ����(#	���0^��]�a�%���A\Yy�=P֣a���;?�� ���y�&w��ٮ��Z��I�2ZO���	W}�C�k"�nT>�,�$1gϚ}/�d��T�G�m��a-q�qvgٹ�I�R����/��¾T�4<I䔮���z�O-����N�cNUu���9�ݹj��U�U���ۆ���HS��%�=�&kz�=�.vٜ{E!6����>yr,��:���lv�ەZ�pb`*�;���.b'�F��ZU�z-O�����o+�z��x�fǙ�����-�b�[X��<�MK�z �������a�7�R�+�bI�k���u�r4zY�Gٔ-��|wMM�(	Un 6�:V�"�0�����~���+	�m>ثW��A'�-�&��J����/&���D����h��8��s.��(�ԍ�f՗���v�Y��wj͜4T���@S���A3�����hH&�x�L������Q���BO�̶@Pge��[������QB�����e�ɸ�` p3TP��9_���VP��V�'�~7�>�О�w+��Q憺P�U�8�O|���jzm�=Ãd
5��lX�PD�a����q��9��:�X4 M[͹����\ֳ��⽡�#���:�+P
~��iB8�t���ȡ�X[��Lw$���Ͻ^q�w{޿��3|]���A� ��C����
A��ލ_7�b��lRYe���2j��ED���)6�5�5EZ�:�K�GC�yK]�I�������I�/f���!(��-〡�Rh8�-�_j_m�d�7Sf[O���/ ��󧰐���ˑ�n�dr�m�N�*l��|8�2o;8<��cLww�KO�$��EG<���	=�`��A�Y��)�?a����7����~a	d�+��`�����Cϸ�up�Vl�D�	}���U�ҝ�Oa���)��$��r-xs��O���5DG��2Ne^'�'ǌ�z)P�uɬ�Q��!����,��	�	�r2���ĥ�p���2YMB�ƪ�R|i�U����,�RV��L����AIVC�d�,�7t+�)y��w���+c�����ϿqE�݋&ҤC���dw�nϷ��q-,�M��i�@/���9+�4r�
�a�*�T����T�?���Ε�{>�]��7~�3>�Q+� �K!h��1ſ�Djެ�<�>�9�/�Z�sV����s��|+��O6��E9Hn����N񙯽�����3�JR�B�׍vWq9IX&����lU��t%�g�����b�)�6<|םQRPI�f@9�v�\��qjZ|D:c�.�677#����Jf��o����`�����W�����nm9a�3�lte��9�-����&�\7�冿u1c��٘�%+T��)c���*�����H��9�Btڞ��"��%��l���d�=�?rTEP[в6�X@1�� ֹʄ
�r�9��k�F�Ƒ���)��t�!P�I[���;�U���P*gҪ����f�u^t�9�<cB(�7WR �^��X�ڂ��Ũ��@�G5E�$ʢt(�h�q�e�Nђ� s+~u_W��Q�&�׼u#*l_�t�����nT������4��9�u� ��ۯ�%������GŰ�� B��8Q#ա[)T���pS��Q�||~\�z�}����(���r<� 6�ۉ_:������uS��N\;ި�B�Ŧ��9�X	��Nf*Η�M��7
����"��cI��(])��lB)�J�*�aq�̶�/M��O��/}�B�;|O��p�=>�ps�L�ف�d���������Q1�����ed\fb���f�~~�P�	��/�#˭�`�������N#K��>�u������~�Z��w��(������p8c�J���}!�	����CM�C����]��2P��D���<#�[wwt�U:R�7_�q�_��U�P���	�@������Y�=y��;Y ��3�������>��&�l��V�l&�c5N�f�p�5�>���M�b[-�&p���O���p~Lkhan�g�k�b���d��c*�/)�H�։6K�e�ek~|���jk��㟘~~�V���� '5��|	f�6��A��8zԜ��/f+ښ?xr�_NÛ��q���·SY[�E�~f������A��|�t�M���O��o-�ϳO+޽��+f~��'/��u=����|_
�5�#���~S��Օ�_\�ԍ��1T.���8�vz+/����鯸P�0�4�J9�#����K ��s�N�����`�8C�pDl_:u/&،��Z�z;uXZ�ڢ����)��Z�r`��{���ë�y��?ָ&ZS������&�M;�&80P�6�+�bx��N�����*��=�a�nQ(Z����[|�����X��l+�~�D��a�P�������ǳ|M���Q��'J�ǫiͫ�*��E#I�=��d)�Ҳf0���OAf�-�����Q���b���g*`�)PIY���������;״	��^���3�Uy�X���=`�l��]a���nb��ύ뚟�]��~l��۶�rRh^AD��۷X߯����֯0G��R�41s��8[n`f�t=7ޒX����9��]�*��3g�c,�D5���L�Tv[��t�~mv"��
��-s�:���5C?pG`�$Ե�oe�[��eX�s�2�O�4��q�SG����*��(��v¸� �f5qS�%i���z�����u���|��s��,;�����g����]���ɱ$1]PG�Cԝ*z>�"��1A��^�Q�K���ʾL%���2NL�;�ޫm-?;ۗ�~�����݊��Ȑ*�#�\���Z�
U�a�N,6qu�t��^�04C�tF��ᾏ�m�6�3�̞��S�%<���B��I;6�����|o���Xt�H47�}t���\B��?�u�?�^��-En�	���mNп�§Ŷ�p��}_^���ebq�����c���}ޥ׷|Z�&7Ko-�����I��?���rQ�f3�l��$E+��ի��6��u2+M���r� �ߪ�jk�Ol��*�����)��Jp�|�-OL��++2���)������Ή����R�X�B��p���o}���I'(��z�z��~�C�΁��͚Q�Ae�^`w+�
31՝Q��m�4ѩ�X2��oǬs��.�ʥ��d�/t&gmbu�阢Ci�+4L}��%�+�����H��(v<�`��*�@��$5f(w�wfD;��a��0%�����3� ��10��+ELq[�&G��sP7�e��m]>���6�,�0jZ躝f.Q�_�o8��ʁ��ֿ��0ҏK�?:���yu���t�@���E�w[WWU&īW�r���u�m]`۶�T��1>�Ms�L��ʅn��.��r7��N���G�n�����tpO{{�	�n�>��6������-gͦ����·��/�p��'&��Ȁ6�����R8��J� ���4�O$�)�#�����Ӡ��+P�O'���}����Ȍ�����X)������-do�����!�6�D���{Db��VlY����$��;�/:;;;??���txs'_N�k��e�C��C9T,U�	��$�޿�x>�-$�Vt��qQ��5��+ri����<�5H�c�������mjj���.���ck�	��U��@J���p������F���g�Za�9ٻ>���Z�Ζ�Q"��/�g�㯵��-RYy��x`
r�i���bZV<�Bjr�,���\��'A@?��|,���ʬݠR���m��!���J�㊬XU�	QĨj{�*U3�E�Ԧ��q,lu2�$4b}mm��V���+��+L(��U]m�>�\�������+�#^u�D
�=b6�.�-�=[��S�KW��*��D)�q��A{����~R/�� �+�p�Q�I[��j'��9i����6��������u]�������J���w5Z�սx,@:����HU-f)6��f�����,L��2-B����k��Pb����ge���0�QO`�L���Q���܋͹R����_�� �ϯ�O�I��M� w׾oց�����B��2�'����#-zoGl
��q�Կ����*M;�z��qt<�5~�n0�4��zn�#e��CO�� ��-���������pn|�ð����~�os�"��]0/�� �����@��IG�-a?�/�zز�}z��q�����t�����=���X���ߡ�.�[�F�,��|L�`�/i�z� ΍͐�W�𝨯�s��@sf���c��6݇��c\�~�qii��Bmcƈ�krTĲy-��	�l]����@�	�qIF��Ћ��!@u�t��-���V�P&�L�?�,�;Sv v���C���������0}g�\w�w@�}��e�7����ݡr�e�DGG�K)�����g;%*���@>_.9���Nb�e�f��Ca�?ۀUJuO2�-�0�ʷ�ܧ_�=�~�=�0~�:u�	K^ujU�Ь[̟Z\$����� G3֋ �9@�p���$����۴6�X`������������;96�٦�zv���I�#5O��߿=^|��3��Ș\]]���0䚷g_���p{~ww'U��_�t���pk]�4�zc��Ro��"��%Jѐӓ�K�[{y~]:Ү3Ҕ<u/��>��;���;�B,i
г7|�\�}�#�7���%�{罸�Ut�/"�Vo�A�<�)�u��o��p���M(��ꬉ��"�0�76!:�"ny�DAfM��)k���}B���F�|�Ťc��#ܓk��������y�h��V�V�unC��bX�m|Xa�<������r!�+5�0��-����v5\����?sl+�΀D��7�If��q�/B���2��ITT��qj�ic��r\%�4qj`�d9{ŮU<h�Y׹#��d��
 �1[�[7��~�`��N�4|V�:�@z�C�%Y���}��HX8^q�����e����8]MR�zv���t�|��{�N$y~��M
"�ܽ�%5ǆvm�t]�&+�
Qs�mQ2AY��d�i��Yå% �Ҳ�IŢ��#�B(�%%�S�A��+�v��˨]G1�Ǣ�n4�ԯ� �������僃�|�'A��q��VV�_�+j'�eR��$H;�����.�י���Q��TC,]�~�5>@d(M-f�5~�&�dY����N�8Ҽ^���7�(!��ٙc�����g]�k�Gn�I�>����Dd�-R;�UAQ����e�ZX���}�ٺ�p^aц؟�
D����	SdU�� �q�6�3f�����g���?jĪP#h���WQ��VP��A�]{ըV��أj���ڛ�{�U��U��/>��{��˕[�s������^D1�潍4�Sk�K��N�-����P϶9����g�HO�/u��✧�8V�S]�"�xF_��J�d��N�2����[[��<�J�n�["�ܔ�&&��s� ��	��W !�Shc~M�1`^�55���<-;ŝQ䣜O���H�v�R�$���!�FH�ٽBH �_�.#�6^��Ir�{꾊p��(����K���7RDu��'L[���puu0{��rG�p�p�e�GA	6FX���o�H�o�a��4��V���N3�o�y�"&.-��K��%/��A�Y5(Bk�0~�w��g��c��Mr{]u{V%�忁*�V��w+���]*���rtD�7�$\��#�p�R���u8;6���0�kN����#��?*�+���؛a��eY��<��&^^��O�T�1+��Mfݩ�UЇ��8�\�2	������W36�.��������C��C�;i�>h��#V*� h��pM������/	-|Ks O��֌cB0��6eQ�!����[A�~��z.��fMe��u���'��t�����m4i�񸟚�Y~!�f�}ˑ����=:�i$��w]Cj�Yv�/�p2P_���)�K��0l)���z�Q�_��(!C1N�����,��2��Z��f]��?���������C2�$�c��DqY#D�J��?�����I�g��N�4!�d��!n~�y`)2R^�h�p��K��W�� �"��U�4V
h���1��'�,Ǥ�Ըhji��3.����gf&�;�eR;� �{zz�,F�"���t[� �d�=lj�
Oo�1 +���щh�%�gݺ�x�˷U3�����4z�N�>�c 9j�(��X%1����>�>�}�-h+�'��������w>�rӨ�=�t�S+ڎ7�+��q�r�����<�Q�ړPG��e�Q϶G��4�������%�{���G���X�{��A�#F��8]�/����z���,���e���-��O�N4b�y�ٔ��X#,Z�F���?��9~���|���Xy9�>1��f����љ���I�o4L�p%��|���Fp_�c��?~]>��dT%�P����?� bџ��SR���a��������@@�!���ֿu�5���T'��}U���6�"T�#=?��E�t.��ag#�xϖG2߃b�i��t̀�"(YQ(�x��wɳ�ȤxO����E�a�p���F�k�/��+c�GVy��{hq��_��|eh!T�*n���$�q�l�5WT����G��tf���淕�ּ���:Y�i�ʹ�([D�i�,��l�Ë���ll�+�ĥ �4v��H��za(@�
�џ���]	W�c|0/���\��]|�~�ɞu���A�fDY~4ڢk��EJ' s��	�	�E�����6�ؙ�;j`�����]=��1D5�&���r4��g�yX+h|��(
m�����d�S,6�h(�,��d}�2���˕�ծ��=���܉2C�鱭7�4�9ґ�76���?��b���ŉ���Ѡ1.��G��p:� s�4	�f��|������8���S�O�0jk@'��T]^�P9�����h����j֛*R{�jh�l[��ef�7	h�Ot%�D���9|ͶF�v��S���T�A'mt��t�?�,�S)�1y�[01Ґ[����G|ץW$ߘS-BL�S��*n�W������$�~Zl�V����o$[��Uy��N1rL�瀌0��_6	Ԧ���T�{f���"�����AT��B�c$���jP-��x���?W��0�q�9꠸;8���4{�squ���&�/�H!�>���)$Nd(�?���	�-�%��9����%�!}-��[��n;����
n�X�g�b-�tX�n3�u�ND�1��\��]"�8'� �$ônK���8���fH�E12û^Rذ����s������xa�z<�9K���U��t�#:w�GP�?����=qJ�v�\nn��ɴs���5\Z��I�3�W���0�i���ܫf/NG�GH��,���b�L傯��"�wA�f-Z7@Rĳy�c}�H���[��?��?s�{��OCk��	x�TZ�l���&�y|�ۋ��j�x����,H����Y�	�m@Έ���j�T� Q��n����+ؠ
=��&�2fI��ԡ,�^Հ;*��Q}JΊ��h�"�S���${;��	��7:G}�B������%0�8�
 KDo%�Nj7���pҁ�0�?Y��q����<�3kI��'��W�;��N�ȶ���N�*���������щ�71��e@�_��� -AU^\䛶)dp����O>B���"�ĳ�{�ĢsT���Cm��5���( ����S33ovZ.G��l$��jNd�[�����k�EX��v7&��n�y�ᑚbR����k\E1XF:�3�%�w'��Cu�(;��1���o����	Y[�m����p>`p�[��#�{�	�0��e��%�[c	A��F?�4��oǮ˵��2-Y��'1I�Q�^_l��?� )��L��藱8�Ub>��P«=x��'l����g8�&LMi���	>$H��Im7��rx
�� 4v;7�N���=�7Ԛ�_1ބ�B��{��Q* �}*�* ǖ�x� R��)!BQJ�^Tsi��D#N4~����{u��wP)!��=H���yO�f��� ��y��G�[Ϸ�%�0�~��i�5r�7��ab���<��'󐾻O9�n+1+������M*R侀���0�W �>
Tii�o6����{z��n)e*Ht��ܜ�q���A$���}�#�8���_U��יu�_���ۖ0�R��0���BŘ���ƍ}���g�����L�'`=�;��z}�§�oLLƍ%��r�a��R���O#'p���� sG�|���(d��11��b$�j���sGL:dm�eE��ʔW�Ɯ��SY[���ǒ��fe�6�\rǟ��a�3f}F<�����V ��m/k���)�t�Yz�|_�	;����Q뒜���}�����������Ik���p�Ջ`oa��%;�&q����@4�}�B���j�����O;�j-��K���\�X����Y�ڸ������jZ�+���gi̎{8�?�٨7��Ѷ��p�&aHJz�q��	��qv�C���2<����H�X�����5�g��V������o�KX�.�,i_6r��2�#a�`ʗ��{D_�s��O4�Om�y0�w'�1r�X%�z�k=�k\p?g�c��򹭮651�r.e�X,\f�=��痵�x~�Z����Ů3J� �sY N/p��S��#��R��Z��|���`;S(���!�X*�/W�Ϯ�}nM	ܖ^w�Y"^'����	�c|�$^)��|��&ID_��Ԕ����F̺;_Ҳ�y���lB$��S��[���L2���M4�X�)3k�?�Դ~��8� �ժ�+�W��6���'��ϧG\�tt�|�,.��:���\�����4�L9wth�U�tGq=6+ ����pE�s�#�$&%mk�����yѯ*�2���&!-e��f!�������#�w���	���ؤ6�sY߰-�����"2agoђj#}��Xt�����nIo�@}Y�X���ǥ!5���UL���@^G�4C�0�c��+дq�Ka�������ή��W���΍we�Y�ȼɔs-? ;d��19�m�|���v
_3��\������D�(#���	b`��?�W���@(����f�(�@��;?��6p�8��2��/�+,�9���
����M�<�b��3w~�Pg'��*���_@�����S���Gr����hO9Q�2�G=���ԲF�������~k���x6	��IN�����f���:iE�����En�բ�yȥ� 8�A���<S\@S2�������A��~����Y[��H �g7���9�Z��{�V���\8N׍���y�W�f��9�1`Iu�������0�H������dp�Z	���?罼{&��q���^K�7�_!��O����T���m����F�U`�d]���nH����[�YɃ�jf¬n�����OM&�œ;g�X��̹N��w�!#��2ql�/�a��m�#,���V�(�+�9�����.�Z��N���c�2��.�6'O�Z����ȑ4	s���I�B���vP�5�X�c\��{5�}�x[m�X�3�!n�p�'��+̼�Ġ$��Ob���Q�Q+�O]�F��B��]�ѓ��0�>��?��^��Ӗ����x��O�>�����tJ�{s�,A(Gt��Q�a�}t*4w�r�N��8C���#�i?(x��k[!zT��_W�u�#-=�j\�f��M�m���~|��4/'Щ��Bd��P0���z$�2z�����o$�w�`��S��:,?-9K���c�tWw}�%�Q��jX����)|��aQ=Y@��J8�Y8�f_Wz�>z�����'H�X�{������y��ְF238g
�٪
~��Nb�ɶ@������(��g��ԩ~T�T<Y�?76660��c+=|3�
̗��>��B"{�������^��m���^}�V0c\��$��+�8���N,��F���f#��Tj=��S�tq<�>��aj�Ou�l9����}Ωl�yG� a��5}I��e_K�DXQ�xd`-�yu�����J��f�Fb�	An\Ү/�)���b�:J��Ĳ0���d?n�QЪZ��3��w��Q����Ӳ�A�[/K�6r8ٖ1+B8�0ғ�%�����B�T&��^���3� !�C̫��lrL���چ����� �0��ܙ�4Y��P5��@ 8ߗA����w��#Hև��xj%��e"�KĨqnY�Tl�d�8����&~v���e�J�U���!��z"lj���������Dooo���^�^__�����8k�R�S��a� ��0�їcb����h�T=-�6�ѽh��3�7~����c(0)y��}B�8	��%�]���Y;-�T��>�����=���I�cggo5N:<c ��折�}7�HI�l���q:�Qw���n����Jt������eX=N�3��9'����J�sٺ�L��K�@RF�x8����9�0_��'���n���}�_�)�1-ҹ������S�o5�ȱ��B������
��rҟ���}�/���f�F�F?b�>j�r��������N���������F��s�)�/��h園�un���c_�{}SDJzz��.�'_��@��kh>r�6!����rw<��V�?� �%����?qSB�.^3/�u��	P.�U|������a�ݕ��#4��>��0����fj�ϟ���.,,����۾��SwÃN7�4��~kk��������јL|��b�{'M[#e��w���}�oww��D^%m�-"$�?����-q=��a�Z���6�ժx����K��#�q!/���@t��敜�(�r�冥 +����)�G�:��d�a��[Ǝ���T-�������}��pK(X?k�&ϞD��T�p�g1�&,�X�%-���<�3�_���?A���y#���h��oأ�y���U{����R��u8�!�W<̽w������y<fyU�_D������l��M'��#Bl�o���a�I6J+C�l��~kh�JC���<I���O�4�W]��ׯ_+2��7U�|��[2}����
��8]\4M4e~�ie���e"|�6�^_ѤVR��!) R�޹��'��:���I�'�1.�80@Eu5>[�L l�I�T&�
��n�U��Y��kX��ڲ1�`=c'�2	���~Y�h ^�Q��~���Lw���E��۠���7�Á"$k�FI��($OtΤ6�P>����B�h�����9����9%�y����3\�*���%��htg~�m���M1\�.��ñ�fw��G*3W%��	k�@K�w���E;�/)���r�3����,v5�@߅7�r��E��bl�Q��;�P�r��\��!�WA��J��_�3��5�K����g̦��廇��ތ)B3�밿q�2|�~\Z(.��id5�A@�f3W���V��q1��kc v�z[t}���K�T�"���}"�����@/]�ڱ�ʞl�>�7��N��,�ZZ[
�ʛ����v�7��¼N�J��K0�h��#������?��Kt�k�Q��0����`#J��ߟ�*	����ě~� a8.u�e��Mʡ&"KJJ��#�Dれ!�J T� �w�b����EaA�P��I�tT�w�x_�迋��*��aOF���Yf��R�-Wwpw�`{����`��/�	Fv�J�[��ݫf_6wd����-���hU}���ěV��ŵf�4�M)Iq������_M(u�|=y���s
�ۋO��� g��}7����A�t!���!DV��`3�+�AF������1u��6y��'��C���z|�V�����"��4J�Հ�Vð���7�~��mJ���<�J�I�Vq�w�I6tp�7�gC��ђf��z���h����~�u:�I���}�D�,i3̧��#�#l闳��T;Aq��ԕ�/�H���L�w�}ۋ͆�����/d�����%~gDm0�.֯ӭH��qiCb�QH���� 2!�Qъ*��;���6�Z7lS3�gT��ev��&���� �K-p�,�ϸBN�`}��;g�m�D���7	߮#�O#�S���+�x�A�����JȻ ��p�Α��3r�B�^�d[d�1������j��7��c�k�wM}��1�r��^�i�v$��}@;�A�1P Y��~�|� /1���3������%�Պ���/H`t�;8??�����ˋ����8}���CY��6u����wn���0��ys$��kس�TX9Q�l湑��%	��n���g/%J���9=$'��`��%z�&�4�.����V<�ʓ�I��Y�ǥ�Bsa4�ef�N�$>��+E�`��:|�?k����1��c=#�Q� %J�W�ԃ��~~����{1ggg�-õ*�Xuup� �b6���Rd7�,`�OH���0`�FƦ�	�Ҡz�-	�\|��O�-Z=���Qt��/;T�'|eb����Wo��`D S���¥��P�.,q����۠�Þ�6������䆍C_��+�B�8�5.����-�����
��~�� ����oT	cNeڹG7��Cȩ����=B;J �ZbG�bC��w�_[Gj���?��;����:b)q��T	��l��r@��7<���B(!�a��'m��B��qp�&@��Ú��'R��iB�..d�/m�@X!��5�`s�L�����CQ�M��0c�O��S!��ţv�FI����H�;(w�{��8|2}�`٨%F	�}p���3����_�jFФT�A���KVx_W 	L_|T�pl�ԸJ�R{�ӎ�O�|�u���o�J��S@F�K"BR�<���ԓrr��ꩌ �" �A'Ɇ$)0QP&fk/Z�������́���S����c�勿�b�7r+�Z>�ʏω,�wK�	��>������D�ۖ_UU�Q8M�Í��m �71w~�Xl7����c&�@P���
?}G��V�΋��R�����)Y�>�I�O,"�����(��o��/{|λf��%����K*�O+@����P4Y"���l>|k4�{���k��/0�+�_��c����辏+��1�dS
�v�te�V>Kb��Mac�M<]�����R����Q��e�c9������t�8;�]�c�9EEEﮇ�A4N ��ь��uw#������+�Oy���oB��e	0��<<�W/"k�a�/^�#a�f��}���o�Zl���|��dq�~6�/�J�M�7����.�?�&?t��������T�>��Qz�H�n#��V�d�0�]��*ݟ�����H�3�y��%6�����A\~pA���Ä�Gأh�%�7L��?M.�\�����}j�ޏ�ms|vh���S�J�|��
�  �Q&Ð���-��������½�P�RF�t>R�0���C� ~a�į_@7�"�8gw�]�������ga���g���*|@e{�;��(N���u�����dӹ��`���Q~Э�3JRO��{"MhB�AA��g���H���c���WJ�<a�}���r�Tw�M��V�_��A6�3�m%:��S��_<����FC����-�m�K;gR��*�����UD�i(�}�y!��q�֣�ƀ�s5ͦ�B���l�����=�3 ��DR�Y+����
��-�e�Y1���ɮ@Ҟ��h�u�08��	��},��TdZ�e1��PSi�)�3?�Q�L�0���<c��E9�#\��Ϸ֏g8����+��! �c_��p~�G���u,F� ���a[�����N�CA�����m�)�R,����=<�ܴM+���ʫ/��]:nb����*L?'�>J"#f�|�V�!߾��tGn��HRU���/���V�����"�o��x�|���9!,d�
.���� 1�[���+}e&T ��e�^ݙ'����^�;�v�c�K�I���맅+��h��mͧC���,]��㕵�MM�q�	��C6^��M�4$a�`��g�^��%mr�Ԕ����IO��2��ս{����P��ֶ45�4d�[<%ee����o���/܇U�e������� ���|��.�2�!��Ytcn"�sq߽��s�4�V���D���}��J �kF�5��<d��ڞ���UG�͓��_{��d&���rࢵڛw�8��+��?jó�PA�}Z��$M]��	�48䩀\��~o����U��Y�M�C�J���Q��n�ǘs����T�0c���&�ۧ�0*5��8�#���b�nnv��I78���T"�D!5пl$��S�R�x�Q�b=6<Q�����ٴy�����P`���@���\��;qåFr(�>8t�E��k�흞ԋO�YtvV�ݿn���@�ϐ',�`�]�OKB�F+���\��p�h�ڳ���p�-��N��uu�gnZPT�|���7�B>
�	0�(�˜���^e��}��`U���&
%#��h2�@q`R�>��-k%5�@�H��b�p,����ǤT�~��I̊�z��t��S(��-�&|j%�4����C�:�|�bg'' ��W<;�14�U ȟ�#�$+:!�t��V���`��)�4�=/m�^tCU-����)�y�"[���ؒ.�N��94xРk��W?����"��7�ů����'��V�u��n鬳�ANā�Jzɳ$�١����0�v맃8k�?]��h!gDR;.^��Ы�r�{Xs��
ŭC�sLu;��K����?8�������ͪW�վ9!���/Ktp��Ocs���Xp9�]6���oWJg��@}�������3�r�"�H��ǧ�ث]����O��Sc�.��-�[%?�5�ڹ��ȝS���ݳ�^��G�HG�N�}�W?�&͛3�{'&&4�
��ȣ!=҇���h��g�MKsss}}}�<ްX
���t��a�Ē��v�p�sQ��+z"ʊ��	){瑍~<�C"�٬�`�a8���ֈ����!똘ӭ�2
�τl����s�Mf����3N�U|�ؐM'��lhp�C��������K�t�F֖��@��64�;�-�K��<}��O�&ؿ描3����j���ͩ[�.��,��+1L���s����=4�Q��WʱP���}���O���m��]��?H��yaDT����Au[x��]�����sZK�o2���f�(�39	���'��{��ei;_hu�g\.�c��GӇ�41�Q�����?��|�l��CΫ�O%��faI#�-t��(�D��RT�X`V��n~�r��8]jZ�a,���TS��I1`��l6��Zt�qv�z�L��f�!SD�5�|���`j�f�Ҳ����WZ��h�����7�͇��i�u�B�B9_	�nn��ܬX��#��:GR��*����|/�6+�2k���mjjjh�w���1�F�*�zn��z��ut}P��ebh����DF�;
@�(���N����x�9Fiq����DX퓶�Q��O<��pI�{�����L~��{kXtw%�Iw��]����N���@G!j�,����� =vb�_7�Q�X���v��0d7֓�)���E��(���J�J����	���QxU84X	�q���q�E�'��%���2%z�"��ov�'�޴�'Zm�p�� ,�?��@�h�����j�gUԺ����5Bx��uo�K�� �e����whK��W���-���sz!��FL��ϑΈɿ+�/���C��E�7
��gm�`^�oDQ��7�NTb��@���̰�z&����V촩������s�}c"RON���>|��K��������.���777iii�$�ωͩ��b�	�ˊS�E�Pm@��������/D;��r5,,�����#��E��w�4|�c�|�	��:X�Â�1� ak�	t|�sy��-^d#o�G|����]�俋�}﫣���i�� ����&�oXRKO�ƢVo����O�s�Ȗ�wQ�j�[���a��s�h~���v$��ll8b�����=��M�b˦�"V��B����ݳJ>�q�'�V8Y@�p�8�7/l��>�
ؒ�~�:#lt;��À�����w�<��8����8ޱ �$v.�>
�t����%�Fm�^=��ȉ6��l��\Κ�Fǌg��O�c���iI��V�I���:��0��WmJ��-�/A+Ff����R�V����g?J`&?>F��1� o/ǎ�&p,|6�����Ha�l���!���٢�\��p�I4�?s��9��Gy@��&�^Y���׬F��8`h����U^��sMuwx���xb�j�SR��L�Щ�F���>Ǣ��q�623sHc�_�! ���Ȓ��|/&����]�	+�ߝn�����%$����@W;���}���n��J�{�,ߵ��a�*�����r0
��_��ݵ����\u�n�3�o���2�]�����ܝm��~{!�  G�����/�Y^p�%����:��|1���-@�L�d�ʪ��u���nҔ�c&;1�<�2`vi��5U*Hy6Fj������h�8�3�>�x�C�_����(�	�U�@�eE��J8� ?�0F*sh�&��s`�K�H�����zJ��FI�� H}����Q~YDMП��q���>�+; o��fp�zP]��O�a�	.����c���(!��UZ$0 Vz�G[1x|��b��I��'x��61"�ȋ�j"�Sa�s�̼�8�i'��*j�o��\ms�ȍw��l��]�o:�c��j1�x�y$�d�`.SN��g�Rq�B<�2{S�/x#Kj&�����e��8�u�U���w���e��/��s��a�=��*�����ua�Y�w��>*���mR#0�;��0�e�} ����J|����N�
s���=�N��r���F?֭Y"��5Y;�NS+U��r�;��cǉ����WY2�����./�ـ�3�U���v�'dQȮ�Ye�(u�Rs�ͩA𯊤벐��1�!���S��":����yϳ�A������wP����^p��_��:� >�v���JGTT�w�e�PeU�0�����@��]��5{��Y�lp┴���S�\3�Xs���d�~^|�7ID����M@@��߿��e����HR��\��n�/ϓa������h�f2�3�'�5b�BdD�m��u),B߯$X͍���Zr�����}�@8|��@U���=t��������X<'"���
ַ���l����p��Є�:�Չ��;2�n:pJ"(�ˇ7�����*�V1~�B68�����*����'iG�[�kE�Q�]��q.�l"q�\�%�$�T��!�1' ��F��i����xIzd����=`�'�Ru_�\�i�[\62�t���uk�IN"�+/(t����2}LA1��[��%�=:�]�_��޶o���r�@��H~ԍ����)u=�@�L���9�fny�;u:,߂e������YG�b���)%5�r��8ΰ�G��3jRt�#y������S�g��D*��4��|7W��.L�_�,/��E����d��"���b�/�V���"���k�/nk^��y1��2֣z�Z����rd����a)�9'�q���;����j8ln�����"�%:��}�g4|��l���֚+e�gz;Mˇ�� }
KM�G�a�����}W�T�������P��=�'��%����b-_��Փl��˦�ł���,B���j���/w�(�:���Q��.�����\$De��Ѭ>_ f��8��@���)Q���S?��~X�l���Q�s-�Kݓ���a�=T�8��e [E�6�&�y�k�j*מd[Y*�I_[Կ2J�!��`d*�>R-�1|���o��7���s*}ʷ�����u���L�c���Cs��<0�©�j0���9�S��k��ٍ����M����]���1j��`�W%���s�Us��yd[7�|�K3/C�f�LFMb.�=��{Ĩ��ƅ��ז�L[�66wGĬj�YQqJ��T���������V�G�fT��R�!���358���(��r�~�P��:i�b����[���Vn�l*�{��읱�8�6��s�*	�)3	��M�I��O�}NW}H���9�Wh0&:"e����ɷ��\XU���z�D�OE\��}���(�,{�q��*�r�!.\����h�a<���)�{���w�S+h�|:�]t�1+++)	�w4�bX�<��8����5\Ũ�4J�3�˝��	'�4p��h�,k�c����cY�yo��*��tv��s���*Kf����/�����İ�)sR��x����}�=C����ΧyO���ڧ��Ŝ�a���S�ڒ�9u�tT�M��������as��ڦCFu'HG��kq2��Ȋ�(�݀�ů��׮Gs�Q�)i�(D�%��������0Bp�\���ϝ}���+��򕎗�2d��Io�^���(��O�J�����������Y�M�����r m�?�I/����,KT,yHp�6�f,�n�Ka~�y��Q?�[�/����(c+|IUL?��o����y������7�]���/o�6Ҿ4�4	L����Q+߆X�1�)�^���[<�|�S����_kg]m~�
�����9�Œ����2��2~�¿*+aœcb]L}vb��̛˗#���`�o���!R�FG�-___cM��DN���~(�
����5)99F�~qK�M�����	��|��g`����dlnm1����]�5u~~>��R1�[Iv`b��(�R�/�r_nk��^�5����t�%�4-������}����n���"ܶ���L¡QicF ��Ne�N�Q�,��'�"=�-Z7�4H�鋜�#Ǌ<�:b����ꑿV��. x��M����ېZCD��h:�O}gax<<�j���P�/R���؍�� f�ًi���@��С6��#r����߃�%f�y 94jU���:t��)���(!�MKhG�K�*�k� 1��~���	�l��Q�w͋�$q������P'GgsEء�N��pU�`�"1�yi`�<��5���sm�G�߾I�E黺��,���І�a^w�=+�َ���&=WҎ�o��(H^S������'��DƧތ���8�{�e�к��65��H����y�9;�˅=�#XD0h�
^���㘺��BO��i�d��d��ܿ�Aܱpk��<�Z�ې���� V�B�4#A���WP[[[郛B�oސ�� �~+��BŪ2G�x��_���O'�`��������hx 3}�t�Ly����ڥ@3u-Eh��w�PR�2�Yuޅx#2���@ Λ4�r�7��O�|�X��@�TӂA�:N��b͔M52���'��_ߋ��w������������ğ�@�`PL��E|�7-����[X�ikҳ�O�H0��&�͇��B͕|���=6.��'ϧ0�-��mw��c{?����e�}���I9�a8kR�5��xb+)�d*��|ͼ X=lYP\ps#sOA<�z��W}��;Џ��)�ah)r]�*?�8��&'���{��C��c�o�Γ�ow�b��q�����	u /�����T�u�<Ʊ`\����L�pH��pY��~�HH}���ۈ*d����N���;y��_��N�r�̪��a���@���C���*M������W4k<J��Z�Ɖt��¹�Y#��PMK��t���%e�vDH���(��V��}?�ۓds�����Txw솟b�l�a��@tX�����L�&�����������\jx�;����[z+Z.�#I����6N�kU��6F���u��굎�I�`ZcI�r7	��*�����^�������j�u�k�rѶ�VOJ̨�}p^�SZ653>���$A]l�o�]ȯ�]���I�n�Z�-f�{c�t�J/av�1&��=��w��J�� ]4�����T����+�k�Q��YJ�O�(�ik�J�Ƨ��m�9Z��G��o���Ī����|[N�o����.��yT-�#�|���$���<�8�y|=��� �{�M3fS���}b">��-P��:7Fn��<��Ow0�;]�;�%Z
�:F�1�g�m�{-�I�6z���op�2L/ KkS%��ϹԠI��pW P�4k#嗀)��0%1���k`g��� �����3���U���(� �xv7���c���Z߭L�Y�qnԙ���U������\-=|�S�$��
��X�����ΥZ��Í�.-xD�m��86�hW�Y���e��;�	�����6�qڿ�,���|�c�BI�a��0�����RZVƛ��c��3]��}��9���&w��|[^��C0`�-�+߸������/r�½�RܾM�Q�gƤ�%�aq�S.J�m}q�K��;c�G��}�΍jW8���P���S}��_P��;��T������*]�w�k���o�]vÄ�;��av�L���.<�V���E�p��Q%~}�P��6{k��jN�����R>5n�����UL7���H![��89��m���ͻ��g�7���ZnZ<�ѧ1ʟ9H��@�]���z��J����R����_$�&��Mmi�}5T�u���|~w;���݁��!��IZ�su�.�euH���̌B����cLr������S	�y�v��Pp���<����:Ь����^�u
��q8�������g����r�@	Z�����QR�|p��C���M�GE�
1;7WT� ��N*S9wԥ�1��P����lg�5h�$N�D+˪j������+���5S�~Mݜw��9��f$�5ƨc߅���o�0(}�����������TI��{�KK.��e͗�r��1��KW��V(�U��ą e�)J5 ��K���3��)R���� �V�~:/����jʎ���)WW%�qT\0�\wW�x���ݷk�N����*��G�-��!����'&�V~O�_٨4ǺY7���̈X�wC�wY_^*�~�^�$D�c&TD�Z�*�H`竂Re|����?��HOO�������Ȭ� q�y�y�ҡs��x���%����\
��}���"H�xIO�ыC�QaEM�O�0,gM'WT=������T{��1�3F��h�z��������(��*�RS�`ǻa���V4�L~՚�����_ ��k�)jwG��p���-!���q��H:����p"
�_��k]Q����+i� >V�]ݗk��<[�Y\n��ʆ]�|B/�y���F3a��'�w�W��P�}^��w}���(�p�5t;>����}w{3T�	��2s	���L����Fr�i�Զv�Y�[ͼf���b���~GmDX����R�?�T�~��8Ѓ�JK�e|�ǷuW�����R�ݲsh�*W%�M9@���-�KV���Q����9�2���`�}�[*�Kڶ��.N��~�GK�ֶ*�7R\������9���(_��3]��*�Si�3|[+����'~�����L�wX�u[�P�s�/�pb��/�Ql���Ia��q��|�i����돊7{�-�K���g�� ,�I�,����~k�d?�|ݪC�s?=Б?��;[͍��Q"����o?"[U�L�!�,nk[�T���!�4�wڮ�B�΁)�h��I�w��φ��O�����,�}��Sl�2�ǈ�RA�qu���f�9�?~�A� !,��~�iΚ���#��J�FIkkkg�ӧ2��|�Mw�ߺ��ʽ��ى݃��ZTQ��M�Q����,���5�
� ŋ�)Rܥh�"-ŋCq.�=P�R4���ݝ�@q�����o`2��$�d�����_�s������Bh�)HK����;rwsڕ��OTZI5���*�@�kc��5�� Rr���"�h�������kk��/;!���la%Pô1/|"����Nc��ʪd�INJ^�2a��Q��̯3�&�T�K�"� ��櫪��wl5�ޗ��E�Q�����=H�p���:Q]��4-���<Y��eI@�nn]h��a|tF^��FPk�ڴ�7�ɴ�����w�7]1��'?B_�0 >DT|�/S֪��ʤ|�PiQG%�0��ڨ'+s�d�UK�X��<ѓ���;��Ils ȑv٣9q2�X���U��8�h�|3�ʩ�~Ԗl@
at�X�%i��'��_�>*���b���^���:W]��o˨���9�|u��I�C���>3��`�^'H��52��kS��[���Iŝz�qvU'S�zWbOPe�m[S�Y���_�Γ �����TAbl*��<*DG�D]��j���d�-`��K �7�}&IQ��Q��Ú�7I�`?�u�eީ��
� ��~�n��ɒ(���O�"���� �Hs��a�Fb$e\_�Rn��m�k*��v�U[4�
";���Ѱ�i���#mw�K�����^p?Z^��C�N��g���M-��$��u�}�)d�=�^�=e�fA<	�G≎���	�h[�x��u�T�$������Ⅹ])�ʵ�u?e)LHq�ǅ@����ʅ��s�zu���D0֣B��VeS������IP��^k$�0⅛�{3� �fB�
ץ|���+��6�)\+�H�#i�B���8����n��#�_�&c�����h��W������?��N��\,�x�^s�����E����{zΆ��a�a��N��}���'��(/N��4�C�����oR�l�О��."`�������v�T�'''�'��C��)��������SGX�f��k�p�Q��^iz�8n�d���+�d/J��l�\ô��4�I����VV}��y��O�ݜ�� ���c"bޑ�r�g�n�_�j�]*<}ga��d8�Qc������4�:槖�=>�-
��~\��B�3��ub]����w���ѿ�R!�}�Y���.�0LC�1�.���ZG%`�қ�5j�6�$T��2�e�%�����%�?%��������M�%)��ϸx@��0(�睌`w>0��8�DK6�/�@�l�n@irB+88�I�DUC��J�$�m�Ć�Z�%���'M��?������Y�7��m����T��t����4̤��#��)ò�x��e�߹9���ئ&RG�ⶫ��,��tm^G��-�������ru96A�X#SW�L�?(Gm��c{?�o��,��c�ꨦZE	|`ȣ+�-�?����uj�:Z{�|���x��j?{�E�Ɇ���-N��N��#�5#�5�64f� {�sL�$�R)�+���B7O5<o�����p���W���&S�T�6{W��C��N$���15|B-���*���O�8���KA�,��z&�q߿���H68I1(����SgY�萄�iد����"bX�E��sF��bF$���&�:�<;E�f�(4���u��.y��x�7�9�>�h�B�^%��P5�gB���8�њ�ݱ�(o&�������,=*z�	�#Zs9>��)����Y��m�\�>�'�Z��}xA�@���[|������c$-�ο�I24�ͣ)#��auEKy�)����-�����'�(��8�x�=<X`I�,���uu$�N����鲾�)����ϳ���������e���+
sb�����3�����+Rwc4���|��z~��c�䋽a�C�����+�M��vKɘsU�'����,�5��c��Դ�`��>��ׯ�=���t�����Q��;�ʔ�<�3����u�!��<nZ����[�h�*C�������ܻ�{����zr��W�i��/���)^J��t�������9��Q������B�Q��rF���P;�i�hq���4v=���W�d��u�lC�&@���x�u�Z��8

?ҹ[�n��<hr�9lMdN�ڃ&d�9�^"$$z��!���s�����:A �+�ɓ{���mT����j� �P���	���������]b)��>{(vE��$s�c���Á���<ĲL*�'�A��_��a5G�(�8�l�F�%��ΰ�dԨd>!�o� �o��}��ސ��`8$IX�'�X�����cĉT�����&2�ƇɊ@#��6^�h�9+�1�/��b�`�4GggV��~�Fgݘg�2T�b���'�p��2	*����.�1cw4�%����h:����T����uK�]��ٗ/_ثuCz~�[`�j���M�?7����/���u�n��͂�y����әhB3�4e{{��m�W�kH�ND$��^�Ѐ��9J�ݼ�?E`5^�"�#�lU�������:D��N�8+f<�"wXm�ιb��2���5"t�WJ\�bE ��,������釧����pH���B��<�0*��,'<J��q���;οr����X��l���l+C=����	S
��h\�V=W�H�(	�
"��X��Cn�ζm�z�L���G��'@�Ѳb�`{�hd�c��0�j��}!��=�5�z�<�5���4�K���:*��!
w��*=F�tћW}(R��]�|���HwI�O���;8C�1F�N���9�4R����g���r��~&Q�
h覼cna�R@Z���B�/����#�(�j��A��h
��p�sNS�7(@^���4���������t��d�.���t%リL����ŉ��� U��Y�Ç�ŋ���IG�����|������3������G`i���k(���8ʷw~yeӖ�=i�o!���
�4a�1��Jt�E�`��<���Dt��"�R��o��H�GA�hIL�!?@�v�������C��<���ښ븉G4�uS}�u=x)�Y!�Cʡr&�b6��̧�E�d���\�xu$褭"��V�-�5"��X���%ƍG]��)���S����n�]�s},�5���k�k�-��˻�6ȕyg6_�8w���Y�����@���_ڬs��z����i�V=�h��6���a	a�R�����������b��d�ͅJL��\�m7�3M��m<�I��Rz���r��)�K��;��A�;UY�7�6A�x���h�QЭ]0A��E[4q�((��%�+IJ9=�	fT��#��y���\Q~T4�Rگ�����:n��@��ѣ��M��/�:=[�v�Q�v�Aq��uM-��qLE�]֣D��O
�_���ox�Y�K�٨%�pԌ��cg_ǣfL1�9�G�3X,m.Ǔn��2>p��v�d!�,��_�+�b�&J��^	�r��W����a���*F�T�$x���=f�Q��QHO�ѿ13��G���<�#2��"����5>������������ܐ8˻;��j��ڰ+�Ґ����ɗ0۷��vGiu�x����T�T�[𹫱���7uO�:n{��3WUvP�a����w���z34������i������q7r_��`�N����	��q$!�g�35��D��Tn/..��Ah�#�\�4���ࣔ��@��常8F���ul�o�{����#�È����{�733Ú����xͮo���Df�J�l��}��x�Cx�S�z:G%�ԙ��؞S,B}V}E�ܥ�� <x�(`�ۧ�J��{FhC��Oqӿ�%v���"� z4;�c���?��\U����R�)	%ϊ�ϐ	�����]	kQq{�eF�p�(��o����1�]f���Ĩ�/��c�H��B�A�d!tP:�bpb���Q\�X��C�s�`�}��d	?�%�T|����4�8�d&aҚ��-�Ue��e�*��W����KKC�t�{慯9���挵�WƲ6�X�D�BP�����S���p�M!�Xi�A�:�+���_+B�*f��J��b�%l3���}LH-�}��G���n�n���M��lh	׻����	d�:i k�U�^��2�t��t��t�8���^%��p�u�͖�����wO7�^ykZ�0�m&�urH~�����l��:.'�i=W�T����֭�H]037y� �r̮d��6�/y���=;3e���o� �EddP0t_U @}�;�}�5��x^�|���Q��ڧ�lOd�ז��g�^�g���ǲ�iW�ncJ��I��Tq}���H5�z.Z��2M�]R2��Ӕ<�nyw�ؒ�p�R=AxE��cn.&z3\�C���Pb�|��wi�a��H@S��B�f=�;��An�jn!��g����dwk_gUt��SS��R��ᕣM�;�8>�Ue�P���l�%ݕ&�������A<#�H:����zE��6TϑmMmҌF˙���y�6|5\z���0�{9���Za���	e����� ΁Q0�)b1ؼ@���UB�.�Mf�+��·�j�äBJJ�H�b��ݿ�75a�O��_���8-��4^�\��
}[��H�Gc�l2~GG���UP!��$C��'g"-���2.��	a�{-�����H�$��^����IDōZڔ��:FU�Ȳ�~n�APb~� �����7��=�b�D�l΂�S�O�S	��]6��Y��}"73�_h���<|�@'�IZ�&�Ga�#��y�#k��ث>�5<�Qo�!�z�������ro���G���vfs����d#KJ�˱d���o�m��| ��p�� ܷ&>�y��LI`s�R2Sф���ǧO']ش~����nq��/�ɧ��������9���!����k{X*����w�e���t��Dǒ�kpp��og�+4�,��jŋ����B�nۑ�ї��/���g���?��`==�L.�e�%Gd�I�a(�$R�ٕ���tyy	���AV��t[;��0�s3,0�X��;�M�m��S�\����E��?~� ���Y�9�z�]-m$�F>����:X��1�yK�)��Q�XD�v�5�TL�[U���`�tl|.����ͷ�e�y�R*�%�YY��*�%���Q�φXw����s���`۰���}B횹��I���$�hG���c-+<&�(�~Y�ӬZV����#g�H
H�r!E�^E�
��tH	�� ��!��\I7����y�$,,�M6�/�r�k!�ɂE%9}1�P�{y6<O��� �0L�>F-�3F�c�<�y�My,d��~rl[���_]�"j��� U�.F�A�r����{�9�����c�4��z���ۘ�RT0BꞞ�$��}~p��8��[j��th��Z�<<<�<9b��P��L�Ge�/�� �Y��+y�^::=�J��*W�\X���|�Z/�{*�����ѽ�dYP	��C��I% �-�T��9DKE��p]~�!�q^��O���L�Eع���urDr��*�������G!
J���-5T�R��KW%K���$�c���ro	LZ����:�u��$ǲ �wRWG�_F� 3W��me���8��w�>���<t�~ �9DlV�Ǭ^κ�>?Ì��gR�Y��.h7h�9?�z�{W5ӝ�XY����������lg�
a�H�^E�%�[�EnXXFP&c����X�cӒ���g}m�z[ ������w���ͭ���kb�������d��[	R�uu'��+"~�I=�//��,��|���j���_
Y�w����SY�->v�c��F������ſ���Uzz3���'��ԙ�3ueS������;;���b8����x_:�J�����+No��rF���³�����Q��k��u��ޟ�B��:�
L�'�?+m���W]}xtE$��_6���`�FD?zymՊPl^^A���)گ85��ΦS�  m�������;޾ձ�A��`%�T6��`� -���u�7G��������x1�kCO_i�"S��P��G6��s|��n���\��I�cA�+N^�4T�W�WN��*2�Q�c$��ԊߑkP\٬�ӱ���|5��08%���dp%j�)$=��D,�S�5����i������}B��5��ឪ�~}��5�E��9T��'��5O����t�8�RR��2�N��),�@���H+$�P��ֻp�Ʃ~��6S�m
.��'.�l�{��G$I�'?��K]�ȳ��kml]9�^ᠧ̞�c�y5<���,��e��ma[U]���mP��v��js�V�.
��,uA���-���?�(\��^��m�%?���� v����}��'�VO/�xV �K���SSP9ͤݜp�zz�{{i�p<����0�d ��$�s}��j��?��H�1<�4.@��%[ZX��br|v�4�����u֞��n���j�r2Gv��W9��g�7��3�1.��p^�.|!�_��X41�%�q;S��)7|C���N(�����q�~W+�������e����ڏ�מ�:�����:/jՐ�ֈg˓z��J�����J�A:�hjn���=����_�s�{aƩ;TFOO����s�Fw7��\	Hڗ/��@$C��
��Fu�Ah��v�����|�0pPe�D�����Cއ��-H�<B����hl5�ܰ@�تp��Жe[�v�kH�ǂÎ�$e\�G{{ܗ�*D�^0�ϒ*�u;��Jt�*>[A��Q�P,��Ӌ����^)d��<]������P��a�aA�e�������yxx{P"x�Ή$+E�h��*��\�U��_���۫`��?'+�W��� yf٢E�UY�ʊ�.^�[i9�%�|�`����0�U3WW��<������g�4���0[�BBQg����φ[��e�ׁ2|O�ܳ�}:��9�" ���QQ2}-��yz��A�[?���(|=��t��=��$k�[�<6f~�|�;����Ȁ���w���� ���u�qe���e."�ޖQ>�m��/��wTdc.�@"ӯ`tlwô�Ț�U��Q�\�Əm���򎛎��Ryf�:�����B��L�?%����nQ��5ygہ���:�mJ�����7-4>Gc�*-KI\
�z59b����>|��D\Ĭ������n<�S��@����^��7&5��x�7�rlZC�OA�3�ئ�(�ߴ�l�S!�~wyx7S���p�0&y1�C q>.q�|��j!BM�,lۗ�D���#�k�f����0n$�5rպ+�)~����_���9;��Q��۩�y�����˺~�*dq���#�i*X������0ޏA�Q+ôҽ�����o�jX8K��+k	�AN6J��n�%A`H�"#0�U����vc�B����
Z��{ee�L�j��/�T0K���՝���4�4�kD�@8yϖ�X#���0�+��w}��4��f=qvf�>��Yz:���/V�Nv��ϗ�#,X0��3�+�T�h�	�̖&�ˉ��qÝV0�,(��p@_�"j7,@�;>N��F�x�MUʖC�nn����ώ���F����� 4�8>r�m��e��- ����zK�B�rK��64m�'�W��̪�8}�"F6 rXU���2u��J2[ɸ�ko��0x��ެ
X����j�;S6Yh���y��c�>|ν�<}A?� �$�V�҅ҹ�����t�3�om��d�CG{c�ͤ�jA147#<�)�X����f	��5A�]/��V�1����1��<���9nAh��]ɴ;H�1�iab���|4%�[���b0<��ݽ����1�j�������Y��Z��)�UU�qT��y���L37w.�����#A���Y���_��݀����@Z��������u�du�87I��<��� b����ĉ�8N?:��i�a
�Ei��]pd�����0�p�f|')�^�<��oM|��v�,�o�n kw��_���y,96�jj�$�o�i����R~Y���M���:A�Z .Ċ�G�:RS��l�������^�m�ȗU*J�
�lC���c[�q�0���q�|�b����)ͧ2�Nj�#>6���=����|	���8��e�q�	,\p`�1*�5J+���]��Ǫ��Wж4�C+V g��(��Ѽ\M�p�yL���&��_���(-$��Wb��z�>vXΏx� �bg>�,)<�J�Jr�sc�m�S��&�����]c�_I"�4��E���ܦ��k�����B}\\\�F��uv���̬,���ExLF��a�j���͉��|ф��;"f��)vi�Q��hܯg	�_���Y��y��~G�\�4"SK���tu�o��qR~��P�gPp��	N���iY���!,,fL�UY�<��Z�i4��#��ǥ1r��[�+�֟�Ƽ�?C��ql���3N����YV��PARQǘ,.�$����a�8+��%�	1a���9X>��������헎�Ǥ����� 뛾N標b4�.w�7lC�����V�7m����������:_������εV�Z���ڱ�'w�o9�k�86�+�(U���������(G��<���ה��/^���-A����71q��S�G�~tz�f%o	�����۟��gh'�~�򇨰O755�^"�#6���qg���"Ǔ��;5���)
��۩oGs�X�؆NY�F��� �i��F�o���j�����y^��܄>��qǠ�c��Lm��o�ƊD��*y(�K����"���Nt��W��ǾF��|���;�����&��]6Z_zZ�|�n�l�{����qG��!�up;J6�-�HtRr��~iFǉ�x�KP?��ϝH�;�*�EQEw�������))\{�M�e��z�IC^4�6T/>F�/H�6**)��8��4���2_9P�+�ֿ��ڪ�ฆ��%P�LY��Ç�-�������2322V W�q~�+G���G''����9����_"|�Jr�bQY������בh�c��73��?:�1� �J��d��#�~������6��!N'�XR(ܨT�rKGn0}��z+$$|�88�Ƿ:ħ�' &�]W.ΪZ���
X&9
�B������je`�30�tvl�,�fU�w���d��=���߿�?n��UU������z����V�?c��g
�a_*E����cÂE��d&���b;�F�Lz�;�'-�#��/���a�����mY���7o� ���)M)�N�z'�5��A��)A�*�QQ�p1t�N�]��q4�;�����)�����%���e�{sӼh�s���%�Y��;� 
�9���������5S
��j��3�7� ���H�Fܘb�����y%��(c�z�;V%�Il�����_#b|�dʝ8�]��X�85݌/���e�*�fK��Wp��,k����ֲ��MWQ���h�V)�o����A��C��j����'/D��)�g;�ub�[[��K��	и ��l>o���ĈV���� ZB� MA:�����n��x%����e
Y��8Et�d��nRX�^`9���;�]���<n�[�c��+~(�+��(4U������d�e�̡7'4�\y�wK�C�F9QwX�e������6����a�Ik���y��b����۫���*����U��	��	��L|՗�k��_o���ؾFYϰ���Y�Lt���J��_;Z�����\�{L�o�W�wO��r��k�p�]�hp�O��@�� y`;9rTί�{������`ɛ/���qD��y��݃� ]���2*j�MbeHi�O#~݉N�pw���x���'����t���0��p��ac+v�b��6J0��<��5&n\D;��"�C��mpM���sYLibi��l�G��j�ɂg�X���7��(�Ӎ%���93�E�J"��ֱ�4n f
/a��,zB�Q���M@�U�J�&�[/3$D{<vVq��U�D)�P��"KDs��	&c�i�*NJ��ki��ܨ���z��u_l�e47]���!6lf֧�QQ�����X��Ҁk��|R~B��T�?Wj�������?	aE���qC�� �|̄w���yg����(Z��\���b����p����3#<�w5_e��C�Tt^��2I�  �N����rPW��mg�����Z�*}Ŧ�0L[zC"6;X*���܀{�����B�&�G�v�H���z�m3_�G���a!%�3��N���ƌr��a��Q߂�oˁ��)+�yܺr�%L�%)a�m���?���nGmW��Ip��I_�����-�����_��$�usǣi#��(���X-�+'��	dX"b[��͠giu��he�FM�DaNd����<=X &���:מ=Z���`�TV������m�Zr<�~�������>���ի��WƩ<Q���\�����<�P�	��Ew�ܢ��Ȝ�E���\�MPUJ{H����{�� �lin͵� ��jbA�y}l�?�mY0k�E*	�M���Vj�c���7�q��+7�a~eHAm��>f:��JjnJ�Y�A�~�ɪ8L���`*L.0�F#O�D�YF��n������ՅZ ��Ty<������HP�jJ_��� B 0͏�6}A��}�`44-�_��r�o�#Xq�y�ȷ"U5]�r��b�v�´���&[̴emsߛ�]��ٙI��Xm�c0��2=�}i�id�oELb2<���eo�W����Y�Q���|Vi��{4T�[8l���^-\�=�(E������C�:���g�l�occ5t��&V�	��p���GIJ��"�	�,ASg_�4�n����R5�3*8Üa�C�l��;6B���x5�)L]2 d�bE�[,�d�:7k-�A��bg�K���A��XU�;�"om����� HCg;�0D�|�˜q5� �/�p�'�f�8I$��ΥG5w��Y��1ݫ�z�Ȳ�]�S�F/��qȗN�v��M���R3��S��PX�C���%?O�c_O"UN�p
�%	'����ZvL�DA�Z�&o����$[O�!OQ��^�`�ꢒ�>K�o�Q㨄(~�B���n� fA�.�WMʺ�89.���(P�Sz~9�T�t�<�2+$��������
�=}:���9Yd�р�[�D	��F�=8T����jWF��1M�Zs��o���I
WV.=".����`����K�J�Ho��������s,���X �L�����⥪�G>.��Y��/�<�kbf=[V���H�KmswD��_�jE��6�)��/����%`ެ�������4�S�1�#H!�7{y��}����M���'x:����d��X}��Cl��׵#���Z�� ����-Ҿ%놌R�lW���u$�ò�{+�g*2ã���Ef.�a�d�>[V�Va��r��I4�I���b�F�0�����~��Be�L?Di�4K�f�8o�9�z�\��(Qm���P�cҊ|�M�����`�#�A���F�D�E�lY�ij��fy�Eb<
!�`�T�|4!�w"ͻ``<R�#��n���%���{80	��	��VGqX��vw#,c;�U��O3�Wi��Yk��������3|�-��7u�1��k}�5sRf�!+�LFs��ց�=*Q��w
�|X�ƫP�������U)�F�a�JZlr"j�5=�[�YYY=_�5�tH§+K�b޾ՠy���
,�'u$S�����7O䓹���{�X�ëp�Ab�K�IA�q��|(�͹� ?&lt�f����Ԅ����֣g�3c��TE��k���%��q�&�p��le䀧��qU*+�D|���X�`���'�"�P��v�[�P{�4����?�k�S����^�{#h�h�?�h����O/j�7��bQ����1��$�%O�a�h'c4&��]N8�:B�R�-�զ�4Tu��z5͎j%���C9u�!f�'�	~�n-Ғ,7�e�/J*��f�;�11�a�vJ˛S&��[��ļ��~�6`K+�3�x<j�/���HR���S��?���5�B�2��� ���1����e�\Ɖ��c���q�4�������Z�~�q�y��O�BAa�Ű�[xc�owk�c�Y7�VxOU� ��SD!g=J�&OD���񞱻s�@φ�Y�VB���s�;-"�ɿ��^�?g2�S5��~���wJ�
_�-o��4UG�Os�q��6��|�@�<�sM�D��K�-羾G��I.f���׌JNӒ?�1�ggѬ��&��8��D
���x�RrEĢy���_*X��e��y�҂%E%�tiiiŉ����?#+�X�Sa���&����S��oQ�O)��ci�^��n6���zgB���ʹu�OW��v�0�:ywd���!�)�tsj�g�^��w�2�V�L��ɴ�O#Q	W��F���)q1=p�022"���N��mf�g�Q��.5Z�5Z%�p˜|�,�mu�D�����!���%>����������(��I�j�����ܧm̀��T��j��(�x�mO�GĶ�rt�����u���������X��f������
���X>��\B�(�׭�UR0��2������?Q;��l*�1��TA�(����z�{m	�F��޺�$� p���2���"D��/�������ܮ�xէ*+������A*!�]ɳ�/����"�`PWD�G@��Мp��*;��'��B��hN��	x���<��A�4���h�JF�5�����ziR��_P`�F����#lB����CP��m���1d�E��w��,%���=Ԯv�X���j�<���GJ�@OϦ��Pv��V�,d����˱m�I�A/�$���R�d+�C�Y|~�� T�W�_��F9��:W_���˚����oi�Rb���""&��Q���������e�޶��U�����4��B�gtR~F0kԼ�R��a�=t}/RI�#q�3��������܎��d��V�!O]���R�����p�ۢ������v�D�)�?$%��Fv��J@�~�x������]������Dr1��r@�{g��R�ijM�T ͭB`
؎�sى�����(��z�w�p&Vدbe�L!����ƪ솾��VO�K��|�.sd'�j�-�Ѽ�v0J{}(y3~G���~J*���L�a��"к-L�����=��!vB�Ƣ([�.���)����i%�חH¯^�3�J�#��L�W�y{����~~�g󋑰�6��a��5�1�=]1�<#�����	�~�Ƥ�6���5ًG��a��=]�1U�1 K��> ��y��q�MYe�7��x��3�9���\��ב�6��	�R���H��?�\�6��Q����I��7PTO�oV�K#�����x�R�3�y����	E�������<�$Φ��yp艒��!�>AiA�~�E����`��wT��g
(^�vo�ʤl�����$���0�칖�=亙}��-��㓫���s 
:��7��J��{���:]����!q6�bS}(�9f��4Z���ޕ(���vծ8	e�:��V�P&��+�K�vqh^��ֈ���6�}q��* ��.���4š�ݜ8�Za�gE������C_�e�J�����b�ξyI ��J�0m����&�H 5t�f�2��!%S�­s�f{��C��8��E��%�SMG04~�]�-�#����^��#��Ջ41����᭵����"/�S���q�F�5R��ˇ 
g,�䫀��G��ߚ�^�}qT�Q����76���4V��X��e�U����<�;�l���Ї���df� �1��i�����A�\5��E\܅��,s���+�I��lXY��\���"����JR�£��/����sstT���=��K^?H��^�neiJ��f��S�Q��`����ύ���S�a[5M�tb3�l�,x����������)���(2�ӐmT��S�X���k��Ǘ��#7����v3L���>�W��h:g[�;9�Kcw��OA*����#���t����n��P�Ŝ2p� 	3�[���$W��N}���Ŝ���I��#�J><Xvص���	�(��c>R��Ra��ʧ�IfB*s �i�<@���|g�S��6ʛ�ψ���H�h�������5׻��K���]v��w.�)M���������J8]�D�,XSr����t�K�C��ڻ�z��< Z�����LS�ї�*Y]���T<�����T�)�+9D����1�@��U�"C��9[��I�D�~V�s���(8B������M\o���T_GD��]�����
� ��9,�Q�q��c�̦��Ǿ��寅�X�]���HQk��'{�ҡ�,E�Ss	�8T���k9�����'��+�ʘ}$W�P���T�*�r�8��c1���C�b��I ��	���x���f��-=1�ʷ�
��gQo'�I��H��2�J@'��փ�U�����|WX����_�����۟�e3�Xe#��6����:@��(�`�l&p����~���0CϦ�D��g}��f&X���Ʀ�'u����P�z�a���wc��ť�BT9#�Hun��T��a�\�> a��Gɳ��A�U���1�σ��bG~����.T��Z��$��Ʋ[Oy׮o��I�����N�<��i�-z�PQ��n�w%����X����^���x�v���5�m�P�X��F�l[�����錷F�d!��������Oې��l�U�0`%:��%d<����r��ާ^R�("B�?�p��?A���
;w̑8x�YE�g����:��G�IM�aͣ��d�1��A��+��d4�����<��)�O����7�%�	O��Y��`�tX%�.�B�-�j��~������$lϡ/�{����~�c���	�f
�Q]�p����sI5�.���24�Z�
J��u�=��Y���ICcFZn4Q`�ɭa%Y�	��P�#Uwp��o�˕�I;]׺��u��㭫�F@hVo,����g�0#9h�� ��h�����,1a�ၝ���P����\<���L�P�u�IS��h� �d-�y'�����&G�}H=�m�����rjx�N��`S4|��!���چ}#i_� ?,�d�S;^��T��6������ׯ����U��E#&�{��"�p�V��=tl'���sc�R�=���<�F���9SȗݮgŜni�>�]J�o���w4�&"LUkL��>��^���6U�� u��S����&h}���,�W�xs����>�Oż��><.wK��~�+�>��:(S�F&��:�d|�by&y���_�5r�$��eNBCy������^e@��hUegU��4k��
�%�.y��aĚ�Ʌq%B��ј>E��R�aO�E��Dラfl���a45��ʍ�nP����k�($�j�ܖ$��+d�Y��s`NJ��l����
}�$������[�"?���O`�-�>,Q5l	+�}�hy%�r��Y����tAK� �T�O$�Q����#9Uo!F�(���??Q3�3'R��؋�O�����������l�V�v ��"�͐ͼ$�k���OL�qQ�՚�r����j�gZ%�2�W�䚐��=U����*�7���Q��7�8K��)�!Z}1��qv�h(٬>4�Y�}�ͅH^�oQV�> ��o4%�?F�7Cq
t�1���f�y��x���&,��p�=m�>ֽ�a���$."$ϓ�?m�}�Cp�Nuh?�L�e���a���#֤��p�������_O[1�kbn�y�n��O� ��e{�� E���>�Ѽ����υ����Us.��j�Ek�?L9?�V�&�
���E����H<^� >����[;���ߡ��$����<�ʀș��}���Y�G1����:�]����y1r�X۔�m��q�m�s+�q�8�c_%��>�eo���gռS��#�����N���W���T�mk��S�؟T�X]��·|.��.�T�t��I�F)
Pd����&?�r!N|��X��\t,�r�Y�d��G�����Ti9���`Yz(f�����J���`>����/)P
���\��z����UG�L�"���f{�0ՊP:�b�Fn��-�+J�D�W���\�Y�۾=Y%�ux���V"��Ӌ#]�,S�"Ȉ)��������͟�#i��+K�Hٺ��������*�!|["�Fx��U���	��G��)S�w�O5oږ�W��w�v��0(Sx	�\X���}�뷻��-�	�v�i/u=��Y�:InQ]R�~�!��!�H��qs���r������[,x�T�b��J��GS������Ws����ʓ�QoE)�
�]~��,��|�[�f����	�C	�
�g���z5Z�߄��9�pC湒�+���e&:1��j��=�b��r�|�b
�4��''����H:i6	,�;�\�p��ʶ�id�K�W��2��{�B.kѹ��klQ/� *�h�sr�p����� T@��$�p��� D���T�q,�`G��]�V����Yqi���'�{��9��Ӧ�i���Os���,�tvuU�.�yn
hi�v*�Pʵ i!��M/�TʩV�a`�������(���n:�W*�օ��Ro�C���(Us���j��zk[[�7��|뭷6�� @� �k{�"�"�F��;�O_}i�̹ᘌ�ܴ��u���M`�n���mm�F�ٓCJE���O?1�%�K�ə�ϟX���L]��MK�c��'�|Ҳ������z��z������\�=qin|�Q�5�*,.[���m��{��f؇�r劈���>��c��}���W���U��F���.{����PR�$̗���w��<�ϯ��cG[�X���H@(C?>�o��8R[Y�=/��V��^j���̕*j���h�乒�,-!A����჏<��V����oZ2���m,�FqY�KE�%JU��a��x׺����H롻vv��'�G# 4 �Hlˮ�k������X��R�T�\���A)�d\���V��[�wΞ�4�`�R 4&�1UGBČ�j���G��oG�R���A��ϯ+5?�����捩K'�,��D�$If!�u�����'���{"�1j��8��8�*��"�n�y�\:{aA��$f��$Pʥ��(���D|��[�|p/#:��R��\�V*�F=��$��s��;Z�'�.k��9gh� �P��N�E�����=��	��ri|jyv���T��kR��u�o?��p��Xg��$	DRix}P��J'e$�~���?|�r^*T��g�K�%/��ٽo����ǮN�%�*BbL	"��L���>����t���o����eGꉇo�Ls%�F���A#H4��ֶ����3����Ѫ���8�S��j 1��?�ؽ��������������nn��RR/W�r�Ci�`�mG��s/�������}�-7������0f (�B%%��F�<��c�����cXN�A�!掛k�߼��C����iBj�(��P� Ą��^	b�է�㑻���� Y!��i�M�oٽ7���bU+�fc�!��*� f���>��λnLe���ʍ�_�H�F�̎��rC�ܙ�� -1�H ��Bi�$I �_z�{o?�p��0��Z=�"�n����Z'/\*� �1�"��@+�#�
!�0��0�]Viy6��e�a �8�RJ))��t��<�h�cB�HA�X�٨W������%Q*�4�Zk!�3./�������w�y��X,B!�A��Zڰ*���[��_�z{��%��"%�2�r9��z*��mG�J��eA�u��y�]޾y��Y� @()�=��tQq����O�"9r��7�02r������wgN��p��������:{���3��O��:�;:���vf2��w�l۹sUo����J�p�wmݱ��7�������'��J�(�_x��Ϟy��㧏�s���J��3q�ڱZ^��ꎻ�Z�ԩ3�(�JC�U;:���n/�Oi�NO��7������s��׮-�v.�fǵ|8�w^�8,�A�Є�Gyd��������Ν��c*S���k����ɟ�p⵷/�}f��blf�6(V|{׭W�}sv�-�������DjJ`���a�'�ߵ87��W^;�o�~��W���{��櫨�;g&U�t�ۚ��΅"���"r�%)Ş�zpۣG7-.̩Ŀxy�Ͽ�ܫg_}�»��ǋqk�c'�ٻnM68yn	:)� 7��%Rp�5jރw����[W���W��ܩ�?���]>se>���J����}�����i��nE�QN	P "hY���'��;*�Z�X|�ع�?w��c���;zql1$c�X�v��W�6�R@*   k �F��':t�m[ʥ���؏~���_<��#�N���<�Eq��x����g/M�D�#�	��cK��J�Z�s�:zd������?��;o�~�ع�O��k��U���eϿu>�-2��RZI��Ï<|������W��k��R�\){c�gϟ��o����2�@��5ԇ�~��с#7oh��XX��
8t��O~b�X��?��G���Ȏb�6=1����=��{��9z��\�������m��x�g���=rw'N��`�R$c����n��ҫ�^?}�c����4�/1��4s�m(J#�F%��4�b�����?����7��+�Ӌ/����[�N\^�Z�#険�3���;���Η|L(!  F@+�! �.�����5kz��R�^=?:}���居�j@��2�R�7߸~����`u}��� �D�J�Q��:����X�k�̗���'�u��|yn��<��w������ �A�!&�I�lV�&D ��.
�X�L����͘n�Z(� @�ZUZ���0N�0�� �:^���k�z���#7m����DH�� )����� �~��\.�;::�m۶��(���cJlo����0��'@�]{wf��o7b������R�b��˶ -�2-SI�MB��¡}�>�����M)%���Υ���1�jN���R�����͵���駅�����hz�҅�����|�3�̴ ȟ�6����Xq�ѳ�ڵ�X�-[6�J�R�z�}��l����Ճ������f���g{�Z#��$Id�/�_�(	w�4�%��uO���d�������N,C� �A ��@��t���9���pzd���=�ڨ��&���W3�z�Z`�������V$!D	������~5��o��w���:��ڙ�_���'�LD�U�����k�TGW� ��g�^?V���}�.<q�T+�$@j��ǏX�T�~����~��r�e(A%����ՙ�ꡁ������Z>1R�R)�(�"� �B�R��?z��V�J�|��o����B���2��������oM����C�����!4�!��P����/<ug�58V�={�k��ř�WggW�f�Ξ�jw���k7��_[�FB%Biša��u�{>���F�����~�ۓ�K�Z�PjT���.��!�e]�MHv�P��ɫ��X0�30�i&7l��Gn�� ?9��o��ڙ�(��؏���J����Rkz�t���N~�Ą���	B�`��sCxс�k?v��充�'/��w_�[)Vʾ�aev�xy����R��[�E��^*b��ƹ��'���@���Ey��G���,�M��7���o��M���r~i��蹑|{Gg�@�{������Gw���|�������w������s�T�_�_�~����J����|���L!^��*����ر�W���}�����Ԥi�JJJ�
�Gn�q��� ������/��׆GǇG�\�z�����%ՖsҮ�ck��3#���)%b���
a���ػ{kw�X8y~�~����W痖���_;y6�tU���w�̸�֒� �0f"h|�#�6�n��k��ҷ��o^>s�����O��4��ϑ6�{�������@J�F#ƑVHx��>~K[�(.��ˍ����_����N�=?v���|!��n�%��o��y���6L4 �����漫�4+,FaU�IW[F��+�eلj��j�����]Da�� �d2�8�}�GJ!l�5��wc+�[g�C��I"�$VZ ��z�/Bh���W�^m�Ѕ��j__Ba� Y[.�{�˲�t�\x��v�'�����ݙ�ly�b~�0F����m[iߋ�x��{��O>y_i��0��������K��r�  �MgL�k���ڃ ���Z��T�����'�=�9���#�3���v篝?svY�HE����ŹYƌ�u�;�����j�^ٱmm�H�o�ur|�pX&憕ʹfu���S#�^@�����q@3z;9�)eGkvc�#���<��so,��iNIK6��ʴepP��O/z�<�߷s}J(�5�����lKv~j��7m��B"����ߞb�#�81L۰-B�ř�^;���j�:�n8�!����ξ�����fykW���Q����/�v�q��t:��4���ԕ��)�b�a϶�6���B(�q��غ�ŁP�p���;]�sN0��B�4^?���뉬k�}Goі��P#����Dh�FK��w���O^		mɺi���R�I$�{�7N�,��ۆ�8��*��5T"�/�e�fk��3o����k�k�]�Y�x�0d�����.L���bwݴ�%l��! ��������C��#%-(^y�ݫ��T�M)��Č:u�sx�    IDAT,��ۧ.��x�b���[7vbH!	���Rh��ޛ��X$���<��r  0��s㥅�^�R�d���8�oKV�rι�׷��=W�UV&G�sOD��~��3W&l����8V�5�jq��S/;Sn$21n�w�w��k3����z��ڶ��a�89:z��]
����w���T�l��-��F�M�K��={l<��X:��_x��h��w�fZ�>�ڰ��葭�&N~��߼��3 e������o���)����-CDF�!"��b�q������Zm~z�O�]cײMˠ؆n4�/���s�Ր��w�F	���a��&�&B���>�S�?�~��ϿwnXK�v�kQ˔�ّ_����Š����ܱ�W�1&�1UBk��H��һ�+S�,����_�u��Qڡ��".�?}��?zm9Lj�sk{��U��7�����@���>_SJ�T��I�\$�oس�4�%J����	�~#`�J���$��BZkB9!��΁�3�R�sÕ!!D�\ p�ڵ$I �(���k�T�*	��̙�w�#lXq)Dn�<���������S�<|��`��)f[�OE�/LF+S�^ٔӏ�y���?ٿc��艆L��@j�ji��c�%���B4%�B�����Lv|�Z�\��H�Z�X�Q1���m� 'B#&������ݝ���T���,//B'��2��zytlP�lXv�1�F��Ug�� c�z��۸ �S6� #j�������酱br�	M��03!�f�I�Xue�P��(I`v��l
1������II0��?	#�������g&E��*�b639�/,N̔���H�w���vu�^#E���߱��Hdx�#Ȳ]��Pn dp05>]�W�LϚ..�&�(������M������S���9����d�29
A*m,�N6jIX�:��R�P�!
�(
an��m���rU&�3�]�I�	�j�,�2-GK���a_�ȋ7v�
 �֒ĀH��d�l����LӔ0�CL[����W�\YTq(�s�P��lӁ4'T����̶������ѕR-$��SlP�f,L@�����J�0����Y�	!J�	 Z3�=Г
�x9_�/
��3nV�1-nY�퐙����*��v�`-�D:t��wp|�b窾��� ù�so_^���(� ���!���'�G���HZW�m�g��(��Y{UwW.�O����`wO:��+�ņk� )�5�N�L=51Qn�atuu���R��כkmE ���D���-��2��._y��47��1�rLfB�ח/\���P�m7�NJ5"@�T�ܽ}�	�ɩW��("�0�8C�0Mn	�8}r8�D�G�w��2!��lZs ��ܵgPӄ���K�g�i�Y�`̰\ȘQ+^{o(����=�\��f�h���a۷�2b�������c�u�`���$TOM��<��[����СՆ��:� ���j�Ygu3X� 7���|��{���[�& H�h�A(
�"�1f��dlס���v`Sv�������i�X$J^�0��-��������|�(� `nnn��ՔR?�a�T(���2��� B 2�"Q|gN�[�;�・�����x�Z���ik��o�uA%�������$��H87����?=V��m"�5�:�c� ʲ���!���R*e2�+����`�*��"Y�f�2�*�j%T�k6���r�$��#)%3xOw?7���/����JcDƔ�������:�h�N9f���a��D"�4�[۔L ��(�i:é�t�\A��JI��֊��eәn�W85�$"�
�V��pH��pb2��N�\h�Bܓm*�1���� �����fWW��3E8� ��$� �\T��3״ �!uҝi��#�!� ��i��-��n�H+Hl�  �p-��"���`�����8�џi����B�JR�t�k����c�L4�9�!5H"��!�2q��\6�Q�86�iUOo�=��
�[�Z"5��R�5�k��� �<ʹ�8�ݝ��&��QClFE�kַ���z�$��k1L%PS�����܀�Ԍ3��ڭ݌ D�(�j:��k���$�(Bjd Ԍ����� �U�$��*LHGϚ�3бl�z�WC*�K����S��tH?��p� �c����,��Ā�X��3,/c���;2`��py�jϪ�:��XC	�)�� �����K�r`6���v����KW��7M��2�vl݂ 3�.���H���(�@k��W��Zc���5���i�qp!�%a<�E�7"%�$%C����;&Ѹ���m��8�^-�����b	"��fJ)�㚫�z�Fhq�\���V#�F:���+��ЃUj��tu�!�PH� �:T��t_o[�U$��ʖA�i)��s	5Ivr��T��δ���
�	
��N�U�롛��~�n1$�qX/��\���������X�@���t&�	")��[6��[�
��O_)�XS�"/
�4A*�dS#���!�.]j�M��I�n��.]���J��'��5���/�C���J��F�r�>sa��4���6w��e, lTg���g �2�r��+?z��X^2&!��G)�
b5BJ�z�.�0M׏�j��ɑ��kM��JS�ڎiY��jځN6�|
y����Q�1����á_��k�%D��/m�c����6�#�rm^)�j�x�%�(6��R�ϙ()%JiM(\^Z�6vR���o(M^�X�3�S:@a޾z�n��fT]ȗJ�q�Q�O$*�e�n���r>1ҭ�}.�iC��iE0�Ъ�*"ӳ}�$\ B����!�a t\���ڴ�ҙͥ8��+c㐁��X��������|Z�D�	PPk٤"�Tպ�b#��w�Z��0�Ĵ��k��d���u����懵�a����R�Rؾ�0I�:R��u��C�T�B����׺k͚��U����f��(�Z&o�I��9N�1"&Oۜ
5��������);�c! �B�CFΚ,"&1���H9�@��7cC��!�*jlٲ���Ū�ĄA �a�$2�X�M+&��۳�c��r�Y�E�6`��lۇ�K:�4&�$1n�JSd�7�ֻ�5�6��k[	)u-��ƺ�M+Z!n�ڲ  ;���4P�Rj�V��i8=]]D+��E��	Y��d�t���;���&��T�A;)aA�
r�NcL�@
�S!��,�쎞~BQb�X�#�j� b��D*igZ[-Jb��@Z�,&%PTnڰ{p�ɋg)�S�*6 �BL�T�q]��Wh뚴�ec�Si�Z܄������m-ٮUCՕi�w��)�f`�%�hl�S�����\[�R���*V��,ӱ���H��\�K+��v˰K��Pk�%Z���i��!�%P*���
o���J��s�.wp�DQ2=�\*׌�6���Lw[.�;�O���)nt���y��C$����I��R2����.^�X.���B!��xaa!��:��	�ZkU)�^�P��˘��P#I��Z�|��`��U��0Î/�"n�����ӯ�[�j�!@�ɓhj- �������Z��~���tn1_��Ò8���1Ұ2mY�ʚ,� �a:���>'h9_������ɡm;w��z�X��6�k:�|"t[[{s�cئ�|?jkk�����C���|5@�r��Z(5�9��Y��aR�Al&��1V�B�=�Z��HK�ťJ��$:l��IA�\�d��B)����0⬭����d�G�[\5��`M
@,X�N��@c���k�M��g5M�_���i�\�8�ˉ�_���]�H�~mq�ۮE1Ð`�!�I�X�:�'u��mㆲ͞�\�2��RzI����0�)D�+���y�#�"�MS&a9P�6FY�7�a���q�V*��2(1�� ��Z�ޡU�(����(I�X "��W��R��0m��ڬ��̮��0Cb�Iq��8�;��=�-@*��J�	1@��D2B++a�8B�l�@.K�M��nq,Ba���juq,Q�Zu��=Jb�	a���r��3	͵gZ-^I���b�`Je�hǉi�$	�Ei�( ��:	�$Y��7a�d�s=��5MRN*eL�ܱT�$I*���E���J�3���4F ��b��u��fw���&v[�c0���mF �~��{{V!C @��c��"N��b	�Vb�X۶6#�jmia��m�%g3�&�h4�Jwf�:	�Q�� %@S�% c�q�Ts[Mu���KO.�:s6%�!/n�H{2iu;L�� ����*O)�)��`e1�j���Ͷr�)�q��D�gp�W��3݅��8��PK�� b(5������"���C	�4e٩�kLIdVHE��-7��m����I�e�!�RK�Y,���T���Q)�Ԋ�!H�  ��R*?�X",�[�l0��X�1�PK�Mvm%*�U"\�j{�j� !�~?���r�1N��Ǐ��+|�G�ib�MӜ��h�!,�8�D)�V�?zyr���,�H��e��eBL��1�8K��\+�(�jP�TKK#B?�·~��BU`!2q|}�v�j��ZSJ�K��JG{np�{x��(�����@_�cm:n{+Ow���*h8tx�Z#�C��#K��8�F$�ll���l�H��v�x����G��P��&� m9U����llcK}m)�( �@k��c��Ņ�J�j�����e�0�wu{W��ӛ3lB9߻wy	PШ^� e�H��b^Q�o��˟���\�WZ��}�`�iֺ����-�Nَ�I�~p���iZ��+�}����{�BiB�16M���� ���G?v�=����u�����Z�ÕЭ-��{W�%b��|qѧ�m �1� (˱�cs5l�a����71�Y ��\&��d��&���5qm���X�,070�Ķ]�q��`*0���d߭{töZ���n�I��[Z�-m�ܮ��*n�595[�C� 1�!B�q�����}��v��{�U�#�3�v2��:-�\�d�+׾���U����B-��(�$�Ȳ,۵���\Ib+��У�uqb��r�L�u am]�6�;׭߼Ν+����Y��  ���ǰ\2j��������*�T�����%�J��==Dѣ7��lEJR���*1l��@�zJ l�..V
 gz���6=e�ӶE�\1����wesٔ�E�xl9"H@���RMBsYׯ�a&a4p`��.�`�H9�JFx[w�������0��|�n�c�5l�����*DZJ�q���өT�n�d2�����l{[�i��۳i!��F!�m�4@S�)�R&3�U�Q���o�,��-�L�����fZ�Y;���K�v�ra�R��%�&Z�HX�O-	g��X�6�ʑᚈ���l&�r�Z�r����H�E�h~a�ШY �q�h	)�� _
!�B���������ⴵ:��N;�\�Ki�X�^��W��D�55W�\w/C��?Z�f˩�L�8I�0���'eb��S]-.MM�L��S����pz>�p5?|e��R�8H���2l�J���L��H����������4#��R�LQJBI��j�.%��ߋ120�BP��G&~�S?}mn�Dc�E�@���eqFܔ�Z<�Cb�d)y�wW��/��zjJ!L`"EQG�����q���Zc�1��bi�ڨT�С�����Y�l������go �+�����������|�O�f�L��,,6���[�Ư�]�|uffF��7�^�0�hy������_�g���W�Ն�2Z��ʗ�x�h}�䥉���}�R�W�gJb�S(N���5�U�c_��o�ta%_�� %��ږ-�>��-եY˵Ο�:^ǌ�JB��'f��ЮÃ����Ef�Z}�/��cۜ����R4=]�^(y����o{��E��'N��H�۠�R��� )%7��X�R�u��[���vw{T�\�zsE���Yğ��6m��i��>5�K�9�MU��2�d�#�u@�RC~����Z�X�����F�����w�!�Wu���<��J	�y*��c��>?^��WXYu�c�_>�]��������K7=r����-�:yi	�4�:�b�i�$�%�;�"�n+�?��|��N��k"������O}��r-� P�佋͘FX$�P2�b�6���H�T}����?��Oݖ�[Z������X�M�_���4�I{�R3,j��'RP��HN�x�*u�؟��C;yub._���TƧvnz��O��gy��^��)C�F�߸42��ͻ���[�YWk�?�����x��İ2�z����_��uH3�D�O6n@�_=u�����&
�r8��u_�����f�ZD�97����]W?��G�<�dlx6�nڲ�^��(l�ۦm]�Z(zH&	X��_z�}i�V� q����%��g���*iBF'j�4��c�1��2M{|l)8l�l���~�Q�idL�e�T
J��r��#�U
y�b�Ss�X�� G������:33�Rq��{>v�nY�1s�~3�ަ<�@��}�Z,d2��\1��u, ��Xf����7m�|�ǹ���ab��3�-���Y;pם7��mΆ'�Ԉh��RB	�����6!@i� �R@�$I�^�H�b��3L�!�@1�mjZ6#���B�X�Vc�!��fGܬcJ)ιi��ϟo4{�0�eYZk�9  �f�gZ[s�ׯ���A���&*J�D	��T�xu����\!�b��"
@8�\�k�^y���߽q����q4�(���z�=����#��g��Ii��l����3;3�Ή��7t��5�=x�#l�X�ݺgǖ#zd�}+c�H��Z�{�^�s�-��s����x�#W��2���;�VuO���Y�q��/-g�|�ȑ��(KA�9۶n��'>�&%�??����3�߶��<���ҋ%D�`J��Y Ng+m�d��Gݜ��r9���Z���G?Z�>-e������9ad0�A�A0�W�m}׬ېs�/>���~SN�V���|K6���4T����~�C-��+dctl��3��{p��o�{�ر״VM�P�s�ަm���8n?t�����#�w��;o���_Ց;���\>;��*t���  �C�	���ZH�n�
��I�mG�c�Vyt�h�-}�C��C��.��߽;|ex�rH��(Uj���,e����2�]�Z*�p���\M���J }�{��{��������^x�˘���j0�0���b�w�S.�Ѧ����4KGxkz�?�{_X;�[�nM9���ر�r6�V*�
�-�b&��XZ�7�K�������ҕ�W�D�n�o<���_�
R���D�������5۶��<���q����/��μ�[{G7v$H��&���Ek�eY�xTR"�4�����$�TR�]J<3U3����#W�&�Ė%��p)k#)qIq'A�@�@���w���hԼ���{��ι�.�|a��ܴeЦ՘�����x�$���������k��uߩd2�_�v��ن�I5M���|����l}�Ƶb{��������ʒ�X&QX ���������vy�MF~��ɞ���~�����ݑ����O޷eM����.OUw����R���s�T��m�6o��O<�qc����޸@��|�����;{��a.�<�L��m3��8�sj���?z��]������N Z��]_��s=�Fi.���z�IM��9��D�e�J��۽�`�Q��ǟZc4�>���ɀ}�?<��W���r2��o�s# ���)��d�K��i6k��5�������x:Ӝ�L�p��xy���#_���DN)h�!�wt, 0�]��RB%��鄛��o�m�s�퍳T��Oy�ǰY�ҕ���;5}�^��3���1�Pb�!����:] H @�Z<B+U���2�b�g�s&��1҈�!��K���B)! !�njM�����>pG7 ��i�x��7CUYðh�*N�  �IDATQ��{v�m�铧\���r��4BN�B0�m`q�i,��r�$C�55m�r�h�1fh:�H��B�*��H�i���_�������~�C׫�̓)��}F�[�D8h�i���ze���.����s��Ç�����O@�����k__�qt�̡���?�oZ��Rz�л.�O�Hu-�Z�� �?{�h���������O~�����8�lִ-�m2�=���m�����٬c�m�@FN�����/M�d*�1/��  ����7�������]h���oJP�{�7�b!E�)i��p��xz��o.n�u���u���w{��E�!�A6���j��u��f{�HzM��0!�B�]�q�3	;u���_�����NzͶ��\rfډd����F����؝�1�����_c���UJ�f]�p��[GtbX&�����j&Ĵ�BW>ɼz����{�-)̬��-�A��.��l�'M�8~��ט��933c�	^��9�z6���w��'#j$��liZ�T!1R�>�5�W����wO�x߅�H'�ɹ�	&��4�Y����t7���C���֤D�Pj`����B�4d��ɪc��ȍ��W_����dja�$�}�1�f�`*����-����G��������-s�F�Z�t��N*c}��?����. D��o�&�$����S���=~���߆��GG�Vh�G�^�̹��a���A�>�W�����������˿ص���������8L=����>w�ҹ����/����Om��hߚ��h}���U�zz���lX�o���_}�w���K?z��}X#@�B�຾���'�eCրa��6"i���Je�0��g��Я�f"���>r����H�]J�$�[i=p�tW�O��k�<ٿf�P+��T����L��On	�ֱ��\��QീD�`M7�����>�K��jp
R7︣=�qe�:Y~����;[K3��Ud^;|��b6��P�[>F fQ�N L�-w�M=���&Ȟmw����K����������������e��?>Wid�v�1�P
(��Y��*��
���j�U�U��i�*6��EI�%RhR�Վ�R� �a]�& ��R����cǎ---���i�" �A�U�iU��N��3Qq~����u��,WJL9��I�t$%���aG1g� �  D���R�R��w�TT�:4JT�`iaq�o`��ȦMgƧ?89�u['��Xk9lC�Vk�c�&�86Aҽ_��ׯ�p�3��/Iƹ��Z��[#k׭��3����W�jz�[�f�:x˂�ZKחk�n��8%2����4�>|��������ӈ
 D�F4C�MM�U}�+X:/{K�au9��^s�Rm~xf���bZ� �\Gʕ��Q)e
��o]�e/���� �JNP����Z��j�2�֏^,8~up��o|�\��_�o��H�R2�㦕0LX��&f���3u�a\��r�:����ʷO^8|�̈��e�0�Q���J �R�d�O\_�o�L_�;������n�9S��U���N~x��1"�L�TZ��/"4MGSr��d2D����S#�iC�y͊�!I�iª�˞���ș���BwWiy�Qo1S��F�t.�+�j˥r��Ժ5i���Nc�D4����<�������]���\W ��^�ݝOg����s��@Oy�a�NÖ�ԫ�����<u���~��F�1<<\�֖ʋBHJiER���n ��Li���F�&-��&��8����]4Ms��{�~v�"�2]=�r�$��V��w���߾����䒠IKa�!�u��LL���{�����/<���{��S�5��?���� �_�v�عy��k�}�m�X�.	�E�Q�x4��8������Ǉ?\z��/~���o\���+���HN)C��i��f�s��=9+�^�N��l>�%�*ׅW	c����w���ʙ��j�qB%�1ez2��p�ښ*5��v��.N��]]�f}1(_4ȑ����>�^Ӓ	+a��&���O�tB�����uyK�j�iheӃ���
���5���{�蕋צ�)�2�f����)�\�n`��Xq�q��\�t�٦��7l�ֻq������4�X8������l:�l�<��	VF��R 8�su�5����-   ��Z0RJ$ W�^�8��4���0[��tpp0��e2�w�y�Z���yB�i��V�0�1���g�EQ �1�X�5�uO��Ȳ���ۛ�w���=ń\U�b�@SN)�<�4���+�(�(��w+�:��Mv���A�h4�����ڑ�ᛶm�fS�Ƌ��N^+�������N_[����������Ⱥs����?i6� ��pvv��j���~�'�-��gϝ�(6�J��|����鋥����q�C��k_��:�����/!�`��(�}���KKKWǗg�c�������wNO_Y���$�Q\���R�\p�Xiv���ox���ݖ��Ϟ�ve�Uvd�O-y���TN��X��z���<���Ǐ{��C?�#��	.b�1ָ�v�gJ��A�@��rs|�9wy����2��ݶӨW(�R)!�,�c�5�!�2kK��7���Km��(�W��8}����<�X�Z�ݘ��Dj:!��a�Y�-�	�t����űڲ�Xo��Ri�-�N����c�#(S�d���"A:�H!%�\^۲,P�ոx�8U�$�nr���t����ؿ�~�إE$��}�_Z*s!$�R �#�X��L��l�_�_hH�s1N:L�D��>wy�����?��j���U���bQC���҈sEA��lH��T�r�貴��6��)�ԫ�������_x�l1�Z:�l4��rYJ�bi�r�7s�[6޺u}����Ud��FC8��p�N_w�<115�O?��O!_z�G���>�4)���k�x`ݭ7�ر�K��|�����
�T�0P��У�����ߜ:seq���|��0����0~ㆆ���~�^۲l�0ǻv�ZۃF�4��q �i�鄗n���7�����D&�N�m���1B�	*�"�L'5����T��\�2�ݲ�j� FS����.|4Ղ��MZ�㸁G�<��H`YV��gKՉ�C��΃��[͠�Fj^�q�z���Ԥe��m~�GƄ3�_��0-0S�/6x�o�0�Z�Z��+��Tk�)�Z��{����b2i'��㺜3 %�Hp&:��U�B��� �_J#��s�i��)���T-�� �f�ẞ�i�T*�JA�}��F���߯뺔R�u�ƘR�����٣iZ�R���RJ�M��PJm�޽{7!�^�k��!��v�U!\��-��㕊����Q¨� �J���c��(R�*�v�m�����ܹ3�L���K�.�J%EI !������������⋋���aDQ��Tf�c��{��>;<<�8������l��h�&�XJ944p�]wuue� gΜ��w�BH�ɕj��|>���BJI��P��` �e���M�
�J	)�b����=����[���O����W����B����u���r�-���G�~�{߫�j�=!DMI�٬�q ��	0�  j����;�ݵZe@J!J��l6�w(ݕ�������iBe���yŊA:��J:]������� `۶��4�c�&��!�RIJ���W��m�P(( H)1�MӴ-��n:�
&��%��f��;��  �X�P����+�9&��D�a�QJUVҕJ%�0!  ��U���i%5B(�L�泆�c�k��z���v�E���Z����Q�������;��i��ѣo�6Q�	�m츴��G7mxP�����v��	!~��W��������@@�ԎǾ���Ā�V��=���.O#��64B�+W��m�<r��~�� ���/:tH�Qy��yq
���C�J�݅dwW²�0�禋����DX2*8u!��sE�в�d2)�����do>ٕ2t���v��h{L�#�� �� TOdgI��2�8�}��ޮt:-��j:˕r���i+Y����:���?�Q�S�;�t:�?0�L&V�ժT*��cC�|�u]�*jq���!�T�9�u]O=]t^lU������
rQ9�Ǳ�c��Օ��5M+�����a�R)��a�U�0�q���;!*��0Ƙ����<!DE�l6������#��R
!�z��R�ҩ!�z�>@�gܩϘ���B���B���;w�ݻwttԲ,e6����raa�ĉ���V�c���ݪ
4M۸q���߿{��l6����E�����ӧ���?77�1B���i��L�8�h�V�=[!��J�R�T2�P�b�5������S�w��0� (;K�AՙJ�r�ҥ�_~�R�(�*1Յ1�d2� (5b���c �(�8�a�0�wΎ(�B,�RWmc������L ���8�fS�Ĳ,%��Ҷ�T*%�TP��*@�8V�#��8V�SJB��J�4]����0�5�!Nc  F�Ǳ�� I'�+�1ƌ1%�g]�C�L)�  �9Y��P�Rù��жm5�S���:���L&yGaE"�w�w/�dl%3 d3�?{����L6-�����č��r P��J��M�6mڴ)�HP�<��o}SJ�� " ��Zr�_x�g6��;�¥�k�L2��(�FGG��t6_��^z釯��+�  %�a�v;�"EѤ�:&:�AE�
����4R�j�0M+�L�W#P2�Tf%�!��jD @ A:ф� �Qi��R�Rl&�QQ ��X�� !�Bb�5�"��z��������X�\cL!�P)+�1�+�
 �ʖ��B���*0Z|�W�b�R��0�h��i�c6��M!�B�2�a�t:��B������(�u�0?K~B���!�k�.�4��Z1�
ܪ�w�j�O$
��M��8V�,:7�Z�g
�RJ��*�*1THU� �!�_����&�DY�!�OOO���BT��qww����  �D"�u�ց�%���R� ��r�X�V��f�q'+\�� ��m۶m�a�y�]�ճ����Q�R����;�%C�1�xdddǎ�T
�1B2Ƣ(R����������q�̯��,+�H(e�N�!L&��s)������8���9�i
!ԯ�@B�L&C	ÐR���86!�eY�s��2���y�����O�i��m���l6)�]]]
3�������R�u��U�M�R�6���1�BPm�Z�iB�Y�wƘz�Pu	B XmJӴ\.'�p]�4M�P�VS��ҞKx�QYvr%Ƙ�	ֈa�AD�ohzDc�)��R��RFQ,t�����u��5k��dV'�S�@�� Q--U�y�����F;����1�^  F|箻����[�����W ��z�����o��S�N �BRJ۶�  �����w7� �,˒*u�S$g,��a �JZ :��R��h�g  ��h��%��0R� �Q)�(�h�f۶Ju]�:ԍʣ��8�qSJ8Bq���9W&B(�k��B���@h%!�4C��04M3cj� PX�4Ͳ,�,�1�	5�v
�
��+)�r�u�N�m��P"��f��iB�sssSSSa*̨FTn�a>�O$
`������ ���o��    IEND�B`�PK   �ZIT 3MZD  o     jsons/user_defined.json��QK�0��J�s[�,�־�`��$C��v��%5Ic���X��1����ܓ��=u@J���54(�&!ymPI�H�$N]���5�|:_����7�G,��=�#�]�F��f�qR�-�>9)yt���{�!��r�D��i���Y�(�H0`3F'�Ș�x�iiu��`��Ύ��n�P�wr�tʕl)�D�����պ�I��(h�Ʈ�{u��<�N����1�^�K��U�`��ć��Aot���R��	e4��Y���B3�b���_Vmy^A��gx�>����|�o�w،��څ=��Vh�����P����PK   �ZITR��j  �M            ��    cirkitFile.jsonPK   �ZITHy"F4 � /           ���  images/6e5c9ab7-aeef-495d-82e2-c4e48423bc54.pngPK   �ZIT 3MZD  o             ��4 jsons/user_defined.jsonPK      �   �5   