PK   'sGT��6  �    cirkitFile.json՝]oٕE�J����=���I��� 3ȋa(��&FMz(�;A����S%�6/�f�Y;v�D���f�6�ι�L��ֻ�~Xw?�O��nrk�������է�M7���]w�w�V�����?O��|���֫��}ަ[6U5[Tʹy��L�v����Y=m7պj���}��4�}����+XX!uf�*��
3DRW��
�k�Q�Եa��B�fa��B��a��B�a��B�a��B�Q�B��@���J�˰D���˰D��̰D���̰D��ͰD���ͰD��ΰD���ΰD>���ΰD���ΰD� 4㵳��ΰD���ΰD���ΰD���ΰD���ΰD���ΰD���ΰD΄������������@L���:^;��"^;��"^;��"^;��"^;��"^;��k�3,�)�3,�)�3,�)�3,�)�/9㵳��ΰD���ΰD���ΰD���ΰD���ΰD��x�Kd�x�Kd�x�Kd�x�Kd�x�Kd
�Q�v����������������H�,^;��"^;��"^;����ׇ�a�}��*����qu���7~"�v��rV�}����~�[�ݪ�����b:����fU�O����橶zv�6��SI���~?JBI}͌}�P:+�����Ni�XN�w�Y\�O�r5�o6wuV��W���^��W��(��t��Y�j�;��X�{X��;��X�|��zײޡt���ֻ�Jg,]��ws�;��X��-X��w(��t�[��-Y�P:c��BF��C,��|~	&�L�d���ţ�p�`����^a�����������I��3��/5�����g0�_$�'��`>���N,��|~a:��<X>����z�?8}�|�y3 �3�?X>������,��|ހ�G��Oq�����G���`>oz�����g0���������3���`�������-R�p�`����.�?8�|�y[��?X>�����H�,��|�
����`>ob�����g0��_���WYїY�����G���`>oy�����g0�7�������3��یa�������Ұp�`����n�?8�|�yS:�_���`>o������g0������g0��0�����g0�_���;=�V84p�h������/`�������:`�������CF`��������Q`�������]X�Z8�|��H�?8�|��0�?8�|�� �?8�|�� #�?8�|���%�?�ۜn7��G��,��|>�
��,��|>���,��|>b��,��|>��o���`>�����`>H���Ͼ�7r���T±3�b�������ӑ��N-���ё���	���ϑ��d�s_5���A�#yyd�<r�\��~�z���_]-R4N>�"(�w]�8�T��FP�o�bm������zbc�?��;�|?=�շ�n��(V��}��Xej�����X�itI����TP�� <�2��U��G������ݯ=��;}����NO���?���/d�P�
5C	�kR3D�P�B5C	��U3D�P�z5C	�kY3D�P��5C	��\3D�P��5C	k`C%���\���a��RVˆ���mX񦔆��!&�~V�)�a�m�	��qJiX�b��x��qJiX�b⎿�p��WX���u�!&��WX���5�!&��WX�����!&��WX������8�����Ұn8��}��}������Ұ�8Ą����Ұ�8Ą����Ұ29Ą����Ұj9Ą����Ұ�9��}'�})�����Ұ�9Ą����Ұ.:Ą����Ұf:t���-V�)�a=u�	��-V�)�a�u��;�ɝ���x��qJiX�b��x��qJiX�b�����Ұ�;Ą��V�/)����{W�'T�u�'��_Q�W�yuഫ�������U�Z.���z����z���8�`-�`g8�B�UA_�������*諂�\��q�kW}U���3�v�㪠�
�r�wƁ�.w\�U�Z��8p������*X˵�N��qU�Wk��<t�	\Ū��1�����	��%J]�إ�=�=/Kz��^�3K�󲤷��%�=�|=/Kz��`�3K�󲤷�&�=��=/Kz��b�T.9�˒�j☄6���󲤷�H&�M�R��,�&�IhS��=/K�Y��2	m*���eIo5�LB�>[���VtFLtJL��*M.�4�LBk���2����\&�5���i���2	�ih�'Q�&�IhMC뽕o5�LBkZ��x��eZ��z���[M.�К��{v5&ir���4��{��V��$����j���\&�5���k�]�(�\Q��jM.�5�LBkZ���x��eZ�������\&�5��J�x��eZ�������\&�5�Ϯ�x��eZ������&�IhMC�D4�jr���4�>E�&�IhMC�]4�jr���4�>�F㭨�L�J��e�&�5�\&�5���x��eZ����#���\&�5��p�x��eZ���,*���\&�5��Ԓx�jr���4�>L�&�IhMC�3�4�jr���4�>�M�&�IhMC�3�4�jr���4�>;O�hʇḣ&���\�jr���4�>�P�&�IhMC�35�jr���4�>[R�&�IhMC�32%��4�LBkZ����V��$������o5�LBk�ю\��¤۱�|#*�ɎT�0�{�ʅ��#U.���ra��H��G�m~��n�kSPf>���O����w�]J��"2���a����ce��wXZ�L<V�ك/-`:V�ه/-:V����U�)����+��K�T��a�� ��0{�?��sM[,���,,z���7��:l�Y���w��}�_�R}�S�*����k/����qu\On�(;~�{�[?��O��O���R�;B	��5D� ���$���B�J�&B	��h!��R�AB�?�F� ���#D�P���Um�lcu۰�M)�!�0LX�6�xSJi�WV�+��R�Ä�pÊ8���H�0au���8�����0q���8V�+��SJi�N�a��x��qJ)�V0LX��:N)�� �	��V�)%�U��q���X��|6
��}��}�����㔒ϰ���:^cu�R�	V�k��SJޣ�1au���8��=�V���SJރ�1q߉s_�cu���8�佢V���SJޛ�1au���8��pة���X����
c��x��qJ�{}0&��&wz��-V�)%�����:�bu�R� �	��3��SJ~�9Ƅ��V�/)��~��O�U�˼U����5uEo�
��`5	kꊾZ�U�j����*諂�$�9wI|-���&a��A_�q��IX�1��ע=q@�j����*諂�$��+��iU�W�IXSW�Ӫ��
V���5��`�I\Z�����oE�K�4��4��4�KBkZ��\�&}IhMC���k��$0	�ih�����&�5��0h��$1	�ih�C�&�IhMC�=%o5�LBkZ��x�IeZ��z���Ă&�IhMC�Jo5�LBkZ��x+:#&:%��e�&�U�\&�5���i���2	�ih��O�&�IhMC�=�o5�LBkZ��x��eZ��z���[M.�К��{]5�jr���4�޳��0I��$�����c���\&�5��Pk���2	�ih�\��jE�劚\VkrY��eZ��zo��[M.�К��gh���2	�ih}V��[M.�К��g>h���2	�ih}v��[M.�К��gpH�m4�LBkZ�%��V��$�����(o5�LBkZ���V��$����5oE�d�V2M.k4����2	�ih}f��[M.�К��gi���2	�ih}���[M.�К��gQi���2	�ih}����V��$�����`o5�LBkZ�q��V��$����Ymo5�LBkZ�9��V��$�����yoES>Dc>4����V��$����Y�o5�LBkZ�ɨ�V��$����ْo5�LBkZ��)�v��eZ����O���\&�5��,�x��eZ��v��&ݎ]�Q�0Mv�ʅ9�#U.L��raV�H�ӭG�\�G=R���*f>��렝��{/-�:V��/-�:V�ك/-`:V�ه/-:V�ً/-�9V���^|i�ʱ2�^|i-ȱ2�^|i�ŏ2y���t}��僂��tQ/W��fsW磁�|5��'�U*_�k�R��Ns�ʧ�̯7���8v������>�cr��L~��O�����������a}�ܾ}���c�����&�Ra(~tx��W"Db�A~^���d�K����v(�����~��?&�|�Dz��<�"����݇�����O��e�{8�!�63~;��;�����D����a��Мu��~�^v���/}C���"�W�E�,��g��X��]_ѐ��+z+}{�ҿϧ�W�̊Y<���$� �J?�\���}�t\ד�ן��͠�����ar��������}�;~��D�F
R�%R�5T�",�����a�ԟ�
R�%R,H�H�	� EX"�'��a�ԟ�R�%R0H�H�	�h�"�'Q>��i@�k��h���ѸF��F9�:j@!�k��<p���ӸF�DG9�zZ�4���s�Q�x�8 �i�ӸFN�G9�zZ�4���
�@=��z��1� PO+���5|<,%�zZ�4��cG"���5PO�>�� �i�Ӹ��8�zZ�4��� ��6@=�k�4���PO�>Z� �3%�4�i�Ӹ��78�z� �4��cs ��6@=�k�8��}���@=�k�����-PO�>>� �B���z��4��-� PO[���5�5� ����qo98�z:�i�1�M�hC��>ސ^qQ��$}��0��D>��(у��AwY�⊭���5s�+zσvM�����̗�b������̗�	�_1�+�|Y>�����_1�+�|Y>���A�_1�+�|Y>��RW�����X>��RW�����X>��RW�����X>����F�x��+0�ф~A&�!J�T��Ť��t�	�&�ai�4M���҉&4��/@�=�S	Lh4�_<M{H'��hB����N'0�ф~�:�!�P`B�	��{�C:���Fz� �E5�S`B�	�с���)0�фޤA{��1�O��9��sJE���hBo��=�s
Lh4�7���9&4�Л�h�M�U��tN�	�&�f0�C:���Fz#�!�S`B�	�	�� ��)0�ф�@H{H���hBo~�=�s
Lh4�7n��Ww�w�9��sJM���hBo��=�s
Lh4�7���9&4���i�M�Mִ�tN�	�&�q�C:���Fzs;�aC���hBo̧=�s
Lh4��=�s
Lh4�D�=�s
Lh4�s�=�;Q�V:�4tNi�M�C4h�M�@h�M��Kh�M�Wh�M�Cc`[:���F���C:���F���C:���F��!�C:���F��$�C:���F��'�C�ko��sJK甖�)0�ф>X����)0�ф>����)0�ф>Ќ���)0�ф>��pF���hB$G{H���hB�G{H��оD8r1�b ���0��Gn_b�}1@u����ӑ�KGn_��g1b��-K�&�w�R/��ptw�p��	�c���o���oM��ݡ�%��
Dw�rѰ�ŴڱE-ZU����
D�j���X�he-א+��U�F��|m��r��k��k1_[��\��̰�_o&e���s��e��y	&�o'^^����Wwϟ�s���y���Q���������V7�o�������n~�̷�|����-*ߢ�-*ߢ�-�.�.?�ϿD}�����w�?�.�)�����"����������X\���C��/h�Mp���������<��q�Ww�Gw�o�����ס|O�7YyS�rSU�T��T�75/75�M��M�����c�ɔ��n���OGw�v�?պ�9<��?u�����H��,OYWY��W�uؿ_��u�������c~�O��v�}v`����[o&?������?��wی6��{�a�����E'�����:���>�}���{\�������a�0�=f��Ꮻ��fu|>������#ƟV���������}��L�T+׷�q�φ��V���|�V�f�����}����E�����%&�r��m��Ӻ�v��m6mg����K����2��=�?x������U�7�}~���j �<�Ͽ����//�ۼ��M{c�L�XVo�yQ}�M���o���\^�[U�}�z�a�x��Β������G���o�����-�~����-��-�~��+���~�Ɩ��o��ߢ�/O��ߤn��M�a���j�-��sY�^o���T��	W��7��`�O�I�&�����^�����߭|�g�W:w�n����V�t��W����W�>��W���W��g��������R���O��������������v�7���v~^1̚7M��g���i�Tu�h��f���nV����
��icӻ�=]���ES��b}Z0�:��`d��۩=qa��Կn�Xs�~U�����p��Dov�~_r�ݯ�PK   'sGT���.Z  $Z  /   images/334a8ce1-1ba1-41dd-b982-9eb2c842088e.png P@���PNG

   IHDR   Z   �   ��F   	pHYs  �  �􊲉    IDATx�̽鏦�u'vι˳�K���lv�����"eQ��ز%Ѷ8�c6< H>$q0@$�'$�̗`<P�� ���L,ّ�P%R�(��5�{UWw���l��s��y�������\���z�y���{�=��
nǟ*�D�����[	   � 
ؾ��� �ԭ����A��X��{[� P��N(�����[:CT o���7A���P Կ9-
�?
7����� ���(7~qKÿ���PAg�	A���� f�k����"  U@UPP�ӣ��8����� ��ٍ_���ʭC�����'�/��gQET ��]z�Fvp�*b�g��!K �̬��13�C `DDD BB Pi����Ȉ(!����?������opިjd�.e��o�� ��p��( �c��N>�L�5eYx�ۑ��� bRt����*�0�hL��9�D �M��l�s���� 4  �����*�r�t��@D"2Ƈ�AD�v��	U4�d�ׯ����k��:� �� �T�x�'�ho,�s�n���(�"���v@5�(*�O�s1F��Xk�DQ1D�Z��>3LA�5�>��>��͉2!�b��n��B���ys����������;��p8�$I!�  �omS1(%ƨjAE������y�EY�,S{S�!�1�
�[�&" ������_���>�򪮽K�1�"���UUD
M��~����/��?��/����s�="B��$4��"" @"K���r�� +"zol�5�2�/�c]�,n�	��׾����]��s�.M3���0p`]��'/|�����~�'���_�|���i�
�H��"E�
D@�J�X�C"�(K�1X�u9i��q62�:k[!*"D�UU���A�s���|�+�N�z��gC(�Zw��@������l~��pgw��NWU�eY���ܼ�$^�c�h�! ��u]ք�ɒ�~?�v��?y�D��c�+�,���G�K��ln\ٺ���=�L�(M�,�T�nj hϡ�JA�&����s��W_}�מ|�I;�h���¡
* ����ٳoݵ�ZF��ɲ�+�y��8���wIjǦ��{��'�y���Ǐ�g��n�mo��.Z����z������dzu��g�y���77�Ӊϻ&O����d���� MG�������˪��}>��~l8n����{���lYAb��F���jqTU��2!S7͵(�<}ߩ���O=V�Wϟ���Q�&����#Aì��@�|������O|�ɟ8����+��������V� x�d$
"!1@����+W4
���˚z�ḉ ����r*��T����Pl�F�8����O~���G�nξ��+k&0�誺�T5b����z$�ν��s��z���O|���|������?z᯾y��Rց����� ��� ͡t҃+�
  <;)�D�[4*[:�'����=���x�����x�������:��	� K���p<�'Dɠs[.|}ow���~�'����w�����/��w��Y������X�" ���
zӪ�mp�LVBe�,*��0�t��悱?��g>y��|�̙�K�!���=}|��X��?��TN�T#�I1����FW�7�w���n��;����f:y�ُ�����rw����޺t!���w���ȓ ��̎U  s;�h�@UA �L����Y0��G?��>�6|��/ڦ<�0���?rt��@��x����P���[��Y�&w//�8�r���/^z����+�����B�v�տ(��G~�S��g�������gp�5�pp�������YD�� 0�Et
�a��g����|&����V�Y�-�<r�cG�{ë�m�2��<�$4�L��4ɻ�4K��ޓ=p��ꙷ߹r}������m��'�~惵�����]�8z��j<ܟ@D�[������"	2" �
kS/w���+IYn�;���{O��{eU�z����WD�!6u]!�
hQM��T���{�zd��{��	���`ljZ�/����W���³O=�ƥs�ߚ�'C�:3�o����ύ�i_����	-� ��Y?�S{����^}ՏǏ�<~ri�����xҔeA�B�Q�Yk `�h�p�n�A������~����X��@W�����'>��������?��%��D&�`�1���>�8ni
 D��!$��*߳z�Ï<[�a0|�#��|��Y�\7�Ա���%4q��Pш1��֠ n4L;�cG�U�Q
"!T�����|�ޓy����<��t=⏯���h�@����� Y��N�w|~ep�����N��
��n�
-�8�JYJUih�Ո�Qc�!6�4����*�U]NwwwG������Ǐt�ղ0uǃ��������w����'<��rK��Ʋd >��w/�q�𓏐�kWE��U�M�A� "���R����],��Y�1��������x<.���u���ȍ1�ǁr��W�#��>%Q�`�n�][c<9�<��_z���p�줆&��h� �J@��*�a��(
ʆ�*�.K|UU��piqyeqшԱ)+�L^�֋/������t@���j�:YX��@���������.'�h8�IRN2�dIlDg�UUEPQAC���**U@��H�������6w�j�
�֯���k�덳�ӹ��vP� ����~'E���YZYY\����0���'UU7!D��H� *" ��e�!k Q��Q��))�JUY�;Y6��}��<:�e.*��k�`�lZ8U �L�5F���J��MYCSZ .XKd���!a�h�U@e&�h�	 Ԩ��dΪ5D�D3��;��\&��枅��n���&�}7�L�8�(9�f���BC*�@@#Q,|���d=�FcgQ�tMn2Ĺn4E�t
eI�1F�kV�� YFPD�=y�'�1ԣ�W)����	B���&��z2�<q��$�7��IB $��non_3h�a6 ;��k�[��h�9#g���=�H��
�L&a<	�I=�hY0 �ħy7�u����1�2q� ���D��	L��"��I��u�k��m�e�lW�9��@ P4H �-�̦�ݹ���`wh�`RM�9:���������4��Ի�덈0�u�fI��6��ZE�`��u'�ƙZ�����%A��9��	� �A�]���`��AP@@#H.��\�J`�5�7��4q��
�z�NF Eg	�*�G0$ `����"�c0εb �5d�GzH8��c,*�Jmԙcl"��Xg�+��"�9E�=! �5V�X�|��
G%g��4䝐5�F�"9��cD#[D�0u@��`M�:�!k-N+;�A���m$
���u"��&i�� �e�bZ�%	(�%@e��0k����PG��Yr��j@  R�jP�afc0M�9��Y�7�4!�9@;�' D�JTEP��Pư7�e�%o����t��V�TT8�PM&í��`�%r`Va�����,A�!L��\�!�sB���XUU�Yq�J҃a�cñT$ ��eY��XEQk���`g8�[]Vc�ج�������Lv67����h����Yc@I�O)]�s��*�95&sy�%�*��Rc�WV��hRU��'D�,�4͈�E�;H��ǆ�&.�7�
�bP���x�=�e��L�@�;y���k�k(��NcY GBq��DEY!��H�Ѩ_�I�o���{kL�&�.�uUTA�Qd�������u1��D��CD�rNPm���`(�H�J��p���}���R��4�LFI����`�WL���Q7M�4׊Ai�^d�	E��U���e77��"�R�XKQ54߳��{o��O(�E�� `���۬w ���6E�b4T�B}q����α�6M�K��Q���g�͒�Y����2V�F4rS�������!j�j&!̯����ƕ�%y�)�3���rn7  ����F8^��~o��B���<�Md��,�bHPTP�@[������b�����e��g��F�X��P��K���=����w�X2
�D�J�){����� �*���*�L���t|q}m%��#Gr �}����Ts�uš�&1UT���\��`��)9���a{D�ݥ��cG�M�/����:t�K���PE���0�(����*� (,�zs0<�����u�h���B9��2:CB�V���TU%%k�K�>K����^�{�����d�$�N�/~���..]-EΈ#4@@Z.��#4�g<���"� ��iE�U�dw`M2�:g�jbPǧIbb��lBC �nj1�#!fy7��&[㽺�M�i�]<v����w�:����.���j�@ET�Z�Pr�dA 4`�EXAD��q��ucÆ�j'�h�X�����*cS�$c�bЦ.�*6}�86�e�$�&�&��Ǝ����W�yg��I�CQx��"TP�ݭo�,J	A@Q ���F�u�>�c�Z�l��b� ��f�IU1G�����gi/���dR�'1�$�%��������'������^�-��M���?h����  � +���*h%XcD�˒�׵�w���7���
	���Ш�w�ŵ�]�$Y\����d<�|}2�)q����AͭQ�l���q�X� b�  hci
T� �N�0����ݴ����gI�h>ϳ�~���ڸB�uh"GD"fx����NF�7�.\��5��5�2uVE5��Q�4c��̜Ճ�Jw�Y���1�6
�jQ����j]K]V[�{�b7MV9�./,�u��~H�q��4˓,s�_:���kg��^�ti{4g�{&jT��U ��!k��vi�f|�vB*�Ji�~0
���
"H�XKH��U��#ֺ>��}m���<�W�WWV��qE]mnnomooo�DA����<"M�&1�gi��2:3�j��Q���, 	�)���%�`�(j�K?���B:�tq~~uq����ݭ����ɓEY�m��MH��dqի��tC��6�'�� P���T���
����%��1P[�!�8 m����$$$E$a$�"��CT�rӅ2�ͽ������^��+���S��Խ��w��α��O?�u�W77}��o��_���eӌʪ̳�`p?�A� @��wޘ6�t`��p� 	P�.T�"*� ��(� DP�:H7�5�K�ǟ���Ǐ=��ٳ�W/g����j�f�׮M�_N?������qQԿ�o�%���sPE 0�9�� r�$9l�e���@d��BfU T4@������}�ɝs������I���]$`���Xg��d4�Y���q�PYbBU�*��*(�^�9A7e�a�!6ˬS�(� ؀!�3S��5��5����N��|o������G���\��nn��X"�N�e��ھfSw��{�N�Hc���U� ��H�
��m��-��18T P#���H�I�@U�����`�I1�W��_�����W_���ՅN�L&#r�q}���k���'H�&�3o���h�3̑,�:�Am]�t#n&D��
QE@А��m�E-Dcp<���C]~���y���B'`g�<y����Ys�����zQ���>W�Y�}*b �R�'�����ه�۽�\�` EQDT@Tj}�(
�
@�L7�q:�޾z��������O|�CO9��g�1�~w0�Mh�p}s������w�����fh����� ��P@UP	�n��j����'ѵ�_f@A#�@D������t48y߱O~��ć����ղ��I,��i��mBE����~�d�˗~慿~�/��ō���&�{�r��yg	��!E�7ص�n`�>ؠq�Z+�`Z&c��*�W�����x����?�����'��Г������p9��ۻ.$	̬�$���$�p����sK����|�3�������+���u���&�����>A�=�7�Pp�oE@l�7d�_U�(#"ss��c����g�N�ھ2nU���v�k{{[�ўJ�(��Ҏs����ŕ<����ˋ'���귞}�C�����ogݮ!,�&I������T��9�w�u �����_FA�l�'u]"hݔ��������Ol<�|�ܻE5����ō�Ky����YY!BKD`@I�*�͝���U��l��MYM���ħ�9r|������y3���$1&Iv#���a��C�A������!De-�z~�_�{N�������|����TG��ի��fr�D~>I�;�E�hQ�ba�z��I����l//ݕw��^��y��{���o�����x��Y -�����:����hm=��x�a�
H��5no����_�����9���.^x���׭�y�䣏�s��\����Eu���m�L���wݽ����ؤ�x�o���NO�6�^9������ȣnn��Y�,�;�;��z�*��,�ժ
���KC����=����w/��8~����r�����k�L,�=��M��]B$P%EF`$�d����#w��]�tu��"�������������������C��m;����
���ૣM��}w�����>��~�7~U����7��͙3ߍa��ӏ?���<5������ABT��yc!p䊥�r�Í<�G?}������{��Nk��>��c��k�B��|�Qo���t��G�a�ܪ�����Ƃj<~����s6��hsq���+�0�y��Ǘ@T@�*+eM���c�YXŦ�N�"�i� �̓��?��c������@�\~�c��Ǟ��i���v,�R ���{�h1@�/�%D"��|�٧77��T[[k���c�=87ߋ�ATaf��1���p��4[�Q��.��8���~??}��x�[Lw����j�O?v��ҍ!p8���p���*�oXH�?�6a��K�;y�ӧN8�!r1F�� ��"0�Ri��c�4u!4u�&w?��<� k9�4�V8���~ P���+6g�|���KŰ�w}0�{��GEd2)�:TM��,(��� Tg��,�����JԦ�E�L&S"����l��̛?���|4ޣ��њ��*FEF�,�����vw6��/�{�T��-Ǔ(R���K�0��DȤJm�
�"(���^D� ��*Tu���(&���o���3�|�x��
  �Q ���( ��\v������{쑺�T�%&�&J�Y��͓FN���ev^)���U!C��4YXZT��+y��]�U�y��!���G��2Y=���07g����$�U�,b�Y#��Ah���Z�q�G`X F��b�!VG�,�D��'N��}�������3D�5�s�A2H��x���Y��&�>yz�7ʐRA����;�3=o��ܤz��i$e��1�J}��;si��g)C�q���������by�}6����Z��:D  B�����7֓˓" 7��g�ODڈ ��0QV1�(�k��4E�H��*DTш����aU�Y�����:��x��$2�~_E�1dpZ���	�yk��*J
���&���&�K��p ��2�!c�I�~Yq�7ߚ�7\Ǉ�-ru�\�m������-TԄ�8� � XDD0Ơ��Ug3����ֵ�U�E����Y" �4qIґ`���x�H�7�n�=�ް[&f~���U��QL�"*��Q�mt]�T �I�iuQP$!L� ���Vр��Y��fh�؀��B�l����o��i�*z��
!�(��U��@X���}�j[�EYX�e����F��)�0�( �@�!4�Q�y}���-���K�Cl�Yd�m-[�D���nd�N+"U����EĆ�"*��i�����s� ��*��:(��A� ���
�AD�R�u��\��Y��
�VD��t��Ӂ�P�'����֜*Z[��I��n���qV86M�#*�aU���X4��vɀ����x n-k    IDATe5Y��Xg�ӒYF������0���l����6���n�TE�Y�s�܅��N�}��w�vw��+�F�yהU���WE5� \�c@al�K`����:ͺ�f  �H�C�8���p��ի�#�Tf&";c�<�p�9r��Ղ�(� f2n��͗�����Ș$2F��z2M�Q]U=��)"#DĨ۵�*M(�j<���KcH�C[vo2�L�U���Ξ�X;��~%�6����i��es�� )	�,��!���W�|�����{Ík�vҔ����c]W (m�ϼ��կ`�km�&���Dӄ4���t4(��A��koוt;���7ࠛ���`��!���"l�,\l�!��f8�^����g���Ho�}1M{�ޢ��w	�0�8�Sg=�A$UD4��*�u�#RU7eوP���Kǣr<��t�7Ν?����U�8p�݁u8��bom�L "tD�ә���~�ۻ{��ţ�"�?�6֦i�O����!`U�Ā�$���QE��:�$ͳn����`w27�[ӗ_zm�W��B9e�Y��sǸa0���-�	` �.//5��<��?�˟��O���g�<[M��ut�9r����1Ɗ�q�zŊ���(D���Yg��om����t4��ϝ���,��TU�M~ǝ���D߬�& �q*<�{݅��~��^\ZZx����dasg���G��Y��8E!�
mN "%$��Q��d�u�E<��ѨVȶ���}��ݽ��]��&Ms�B[���Ί�v[�{D�d�m���"u��45���[�掟8����/^؝��Y\^�U�x
!@�n�;�X�Z�Ɠ���B$
�Y�e��6._ޑ�����׾��W�����#�5X4�l���5��O����p�(6J��5�n���p8N�,������㥏|���^�P_�����,�����O\"!TU��ު V���aݝ_0&�ܞn\]���--�\_�}�{oO'�ࣀ����j�����m��
Y�-���ι�.E�"M��K�ʹ�����񹅥�.&W�7���*K=bZ�SBeU�I�;��fgsb3UEa��)'/}�W���`�0&�&S1�DhlKq!"k�%4��ҡ��?+�`�4�!������ym�����c����ǎ]���tzݪ��J�{T"'iJ�GU�d���c3ؼ�q���&�x���ֵ����=UFDDì�R��ڶ�"C���}O\+�QU�$D�֒!� tv�·��z������?�0�_\�����=����^_/�]�w�����3g^z齋�b#���6�tS���Y�1H�;AZW�!�~��:c�����������ΖU������Ҽ!��=�:ڼ����^���N-,�?����T`{{���F�����;E��OTj�pM�RC�,э*��q��p�X�t�}�WTU����\��y�>p�#=����kUYHp/���F��'ww�駟6�>��'��ɵ��ׯlGC�hHXT�9(u�0k�&7r������7�m!�CD�
�L�,**�XD��&�yQM�{��}���������<K�򕯎�#c->HY�}��[g�������׼K�����U�HU�����B kma�T;Qw�9x�[�YP�"GFX�::�4e�M�j29����O�ud��/�������|���'�	G��
A���<��O���N�Sk�1ȑC� �TIT1�/Xa��ɲ_�@���A�	Z$*�(E�������v]��aqy�?��t��-�,*:�ȑ��w�n/'C�+�֚�d�$�*�P�4�ќA��pw*��vX8[�-��}��"(��DE��(�m]��:�o���x:LF;���`g<a7�x�ϯ�/C���EQ��]iB��2��! ��b��~��<���JAu��/�����oAU@�&Ĺ�E��}��ۿ������[i����&!.-.mo�n]�~}�yt�ȗ������Ν����,K"�$�Ϯ1Q���9�>x}n��B�[�B$��R%$BmKǁ1n0Vq�vr�����`)�u�<���%�±��H�Pmv�_����瀈l�f�����B�$��@������[	wFI���v�����HD*�H
�trk:K��>��C�?r���HZ����b5-8�i�\_��}q��3g_~��K����~.�6-��}��dH~�P�3z���PTl��)�h�g��L`�Ҕ�:z�����{�y���/��������`00{��d<���x���}�ć~�s���E��_}�/��W�=?���I&Qbd笵X�M�����2�s�v��R�VAB[�H�*!��/�	���/���>��O����֮�����cE���LF :,&@�W�6����S�������O=��O~����K�����BQ��KT4���u��i�g�QAD9M]�g ���}����e��~�����b�
�����b@�Ө=��C���_x�cOlM6���������,ϫPOdˠmR����R�!G�����/��랇�}���ԃ=��_�?��D��ե���0���彽�$�]�%
�-�Oi��X�������hM�zkw������'��~C����đq�wd����kƛ��k!�DHdR���O-_޼�B��Z�k�~��^�˿��W.�z����t���,A��=��'vG,Z���}8 �A���8�{��O}�g�W�s�ʹB��h�g�I:y��G�� �	F�;g�5����Ť��u5�M��xz�؉���'~�SY7�������SJ��8g�7�~�&;n������m~5VMA�����|�՗!��U���_,�b,�0�D�h��Ȧ��Q���|3��E鄂_����hZ�\=����9 ��/~��������h�:gڳ��0�&;Z ������QAUA���~�9�������սz<��ú*��T	;�3������ 16����u���aw8��4U����8L/_���?x������/��,K%r��`�5��rp`�}��ap��?"��>K��'_8z����f2׹�uu*M:ם�ezg��b.C�9Lʢl�:4uh��4�bp�*�M��:�Kk�Q,7���݂K�M>��O�����Á��ޚ!^߶��~�H[�t2�r2T�&��@��O<��Ǟ�Fդ����BC���-,/..u:=�.�6!QQ��!�X���]�#Έ�l��_]�4l����x\O��xqu��_��OS��ێ���^ct8n�-'���K��}��?���&C�x1jrk3o�e]g�(f!� �(��Bf���<e)�)��殓S�k	㲬�������?����U[a_�ڷ��������I��Lpkm਄s�m�/k�&u�;V�b,���VeY�M�G� ʢ�X��U�M�&*�uif���i��3�o�M�Uu<��S��-�!R�U��޸{*�h�m���✀(�奈R5MY5E�eYTU݄�A��a�1J4(�(�
!�*g�nwie��?77�N������/��Ma�"r���'����(玬��N��>�]�e�q��EQ�؈֑�(u[Y��VFo��jD#25 MC�V�'����M{�Ww�zWW�W���K��錬���;��'e����=�����B8��Nf�OG��$DiXb$+H) �H�""D�$�*ai���14QD�wY���u����t{�~�u܏zo��6���Q��D�����G��v�y���QUL���ib���*D5�0�2 � ��*,���
�* 9�P�M����u�&8�VVV����KkM٘Y"��P��p��8�A�QQȨ����0��3i�ַ�GE�����U0(�h�1����u;3�"p���ʍ���m�BS����H�u�����n�*�iF�m�����SD�7L�Q�zR����4��v�6����F6�8gHP�؀�Q� mA 4�-&�л��3T�$����u� *�1��<IGc�,�*�_�|��rHO:����
Xg���94���'��Y��@BR�u��Vu���YaE@�Dd�C�y��zrd<!qd�QPBS*��1�a�%�*� ���n��QQTh����O|��&*�*1&��w{���VM]��aRM˪� ,���\�$�\7��$�΂����E�ؔ�������("*
V�Y�H����0�"�QU�����0c�e.A���9�Y7�S0` Xߕ���c� h\N[�ғ�}�'y�5.��7�� 
�@�%�O�����6ӌ��� ! �&
H�4Ŵfｩjum�La�B�d�:kcI�����Q�R�6565����D� �`�Q�&d�U��
 i�F�[�r3����1�"���"��r0�&$��ڠ�#cc�#�X��cQ�>K��%:c,�T�D�(4	�UC�(�ZB�F�a��f��os9T������Ѧiʲ�����d,`�4̬m!���/P��N��+����8"�֐" ��b#ޛ��Ԧ��X�t8���9�`�px��r0�`�<�h��X�~�w��w���� f.I���M�u�!�V1���p2�q1�C�%UUEPɻ@m]��A��z.�^ޱ@���<�&�x����V�,���U��r��+E@�, ���6U�����[o=���� J"���ɸ(
�v���R���h�7TM% Q9r$�2$�@{6�`�k,T�3Rg�^�1�����$�
��+7���ͥ�[5,�c$"���l�ݭ��x��{Ou�)�Z��vʦ)��
�LM�8�N�Ŵ�Z@�� �3jU��Y��'Bh��`�߱dv�������q?��:ެ��x�{yG�"3��!"L���������+kw���>)����>ݞ�&eQ���kKI� Q��8�`QT���Xj��n�v�O�O�O��le~q����o|k���$F��D��W��9":(7��p�k븱 ���ޗ>�Y^w�g}��߾�Jݭn!	5XbXll��M�C�d*3�J2��? U���)����J�8���I�\�c��I�ev0H��j�z{�ۻ=˙ϽW-!0 $;3s>�n_u����<��,�C)�ZcΟ?z�=�V	��iZ�XA) Zm8�A�����i�	a ���{q�RE���\��Fi�8�7�8z�_~d3�¤�A޺�"Jc�1�]_7  cRHJ(g��,JiԊN{+(�����+��Ҫ�2OHB�r&B(�U���R A���Y(��DJ,"a�KA	թj�����Ͻp����a����@Jc��{G?��Pj�N8R��1�<iL�07�r�l|Ϯ�RYY��0�Y��Z��j��(c�*��Eʸ �	ϣ�KF�
!�	��R���t��W^}�����6S.WZ��0Ѿ��[k��,Q�
�4�N-h�p�ٜ=1�xH�۾sr�X��Tp��4C�I�0h�X��"p�=��oH���痥*k;�l�3�։7^���h��
8f��%���R�@����B>�e���}��l5SOHJ|���]:����(��}�����F�{��Xf4���ZK,2Kf1@[�$���h��Vμy��ѷu#��%�QR� Ў2ƥ%��������$I*�D4=d�k���=::*=O��R��f�1ƬE���Iñ��y6������=S�r.�Q:NT�j�F+�~>d������L2V�r�<0P(��h��܉��ξu*k��L�aహ(CD��1�|��m�1�e-^?v ��6�/�ر���8��B�$J,"�q �&S+��Jg�7޼�:P-��v�r����f���b*8'�R��A�\��E?��Lԩ7N>��?Y<;2��>&��� %�!@<�K�tdd��1�8s�>�*E�����������y�\*I.Ҹ�qn�5�VJ΅�IV�_\��K��jY���������K�Q´v�4�8f�a��'ϟ�=s����@�	�h�j]k�k�!��ɵ����߾}�v;��eY&��~�  �"����Ν>m�UY�����QGJa��R�)���~�e�K�o�jG������`���F�X,#�E�J�5s�I.�LG����$�A^x�,j#Cp6��HE�j�S���f]M�퇞�@�5� ��_����f���4�(�Z)N�����<dI!,伐+({y�t��,�������n-9"�&�*�P�ֶ�"90��"8/	qm�M�T��~���� ���j�ү�܅�������ɓ�++�g�Q֢�Rkm��'ÀK��,�I�hQ�������[�NdJ�J�]8o�5ZK��j�#��\�60�^o?~l���Fq�u�@!�1�r�c1�л�������%�4�C� `_��W? .!7n��ixd�왳K��B��e��{���RH>�b�w��W�������S��u��ˋ�gN���$JF�~�_�}�m?�������z}=m'� L�60`���$DX�X��g?�|�T,	!ܚ�֜��_͙P���{=�}����K/66�|>3�j}�k  |�"ęs�r�Bmp�ӟ���ӧkՁr��s�4 ��S��j�r��''�&F"��,��mk7�*K777�QښNԩ<v�g��¯<�裔	�,��w|u��U�SB��R.?��SSǎ{���?}�T'�l�o���������Rx��`���ml��q�v���uJi���@a��[�B�������Ή(ꄹprǎ�ff�y���[@J9�ң��sjD����EJ��7��sî=�~�ӧO��,��괣'������s�;I�r��~z�G��T*�\��/ln4���`����?��?�Ϟ��>Cb	%O���}�s�%I�r���+�j���Qk-p%����E������Z�5c�1f���,��������[���_���|���Q�?24���<2<R(6�׳4��X����eW�a� Q�K���?�����)�!�y��ZDtB�˜_U6���] �@��Dp���(#�!�*���>��'O�5������/dIzt�h�P$���B�f+٪��h��T����fbrǓ_����X�u$����"S�-=�@�cˢ��z|`�:p_��U θ�"sN�J�I�\R�}/�ٻ�Q�	/IS�(eC�aθV�$�1��3��������ؾ�J�r����Մ� �|��v�~UT7D�a�*�cK�� �! ���% �SJ�D�8J|!S!�$� ���:�JS�13�'�R$�$	c�x����(��&\� �^�R��5�p5����/����*�)R��j$�tZW^'�@D��R�@J,�%@�.����<kL�ӡ�rƉ%�r֝�͗���p�t��_?��"�ۺ��!�L�� n�&!�<#����!}�h�W�-�a���t���^�V���p�/�u?�wG�V9"�����;`���,��KG�[�����-���Q:\�e=����}�]�����k�3o�v��}�GDc�Rj��͋��p�R"�����qE�#�����']?v������#�������jh��!�����ޥ�Bq�!�kJ�I:zn�Ͽ�tM������F%�\2n���pƯ�w���ܭ}�ݫ��^�ʯ�*E�Eh�՟�.$n��Ͼ& |Բv��aL�e�C���]Cvl�J)�/�=\����]#���qE��e��|���~�t��[�b�QZ[ĭ���x?t���E7�8~�P`O�^�����I0D���)l� �����8���~������N�!!=#�c�8v߻������#pÝ\��b�Zӵ�,���^ORW_��'�1Fc���]�F>4]�3�E�yii�{�����XB���sB)�h�{�;]����祱���^+��,�x}6�5������g/a�{<�k1�S���O��5g�e��ʩ��kJP`́�<M��zd�c�c���y�Vco�t��`Y�M��j���
�"�(Ƹ��>[B@kݗ!D����O,�\�yƥR�"L���a�����:�9�d�Sp�Z�G�F���H����e��. �~���>�|O���Z��.4����4������ȭ]���ԭ���<Ls  �+��IDAT�_�,�\�c,��\:�~-��Lr�����l}��
!�VZ+��9�q�:����l�1F)��1�]��1�-�s�&�[����,=@�)B)��s���~+����b.GVBc4��]�eҍ1� 8"��Ƣ��R���?��~���q�j��f�w�s烼���-$^ZZZ\\�4F��H�1��RD�� �ڋ�v]w� Zm	u�(�ǐ�^�eo�vPJ)�JřN|�EC��>V.s���k蹌�gs�
��(� ��j���+�Νs���P��NvXk=O��cǾ��o}���T*��@��)�k��yN)��XH)��3�z=6��jmA��q��-�R{�}�[_�֙�ړ��Ie�[4����Fc}}��ngY��6ZkmI�$�/#��/[��1��l�ɡ�'�di��r������`\e LLL�r�-���n״�m�ua2ƌQ0�K��B9P���e����������  �����x�[_�Dkm�i-�`Ld*9v���Ç_{������v��6[WQݪ;�uM% �=V뫂I)���Щk��bŋE���< �R�A�sMd��+e�	_0΅Sn�qϓaA��~�Xܶm�޽{o��Zm�{9��{��2�]�M���g�y������c�677�mf��G5�Z�}��v2!��RJ	!�I�(���"H�K¥�J���ʔR�������rmL�$kJ��"!Dk�� �ec�B�X,V*�'�?��O<x��D��.s6��\"I�,)�gΞ�����7�񍵵�j�*�t�-cƘ$M�� �\:��5㶃��R��=4`��k��2�����nt}��b��ra$`}Ngo�SJ�R� �Zs��������Ю�{GFF;�����t Z_z��~�O���~���a��ƽ�v+���r9�]�����j6���h�U��v#_�Z)xf�a(���,8t}����X^�*�RH�`
)8n��1VM% �2 I�Z���1�)!�b�PPJ��M��V�q���f;�#<o`��9�]^޾�����R�>u����u���c�� ���}����߱s��R��e�1v���S���#Gޤ�v� &�PYF� ��(�D�4J �`)bjĸ� @� �B�(C����d�+�8a6�	�L.��$� @�6P(�'&&�����ΞVfF�97���6>611^�	! �Z7��M���ELJ�����}�СC�J�Ӊ<���'?{��wLO�,�ˌ1�������]�����<�/��gϞi6�B)D}m�I�cpO|�;��ps%�%�  釁(�%�r��L#1�����v��{Ͻ?��[o�m�6�����걣�^x��=���'Nt:������;��#ƚ,Ӟ�H7� �����m6Bȑï���V�P���~���Ɂ�j�\qz�ʘ��,�+�S�SS�q����mw:�fY��uM/@w6�)�W~�+*T	 !����XDK��p!��ʨRY>_x��G���/?��'&'&˕j._�RT���s�M7�s�4���ϝ={�V��߿?��W�&R �=vٌÇ_����b�^_{����o<Y(�$q2���Ec�������s�ԩ��~;�2Oʋ�]�[?�O�Z��
��k�" 8�#�@Ќ��|�3���~o�]���) H�7�dZs!FF�}�S�*������/��ƛgΜ��Rhm��ww����fc���l��X^^޽��x�P(�q�/���m2�X�	�V����q�wnnl^X�@�����PBqKQ~(L�;3�9w�6�$N�7�9�S����|�7s�ݭfCJ)=/�"�R!F)Zk�ڶ}�å҉S'�x�ͳgϬ�� �4��9	vw엇Ӎ�ͥ�%��e�[n	�\����he���K\ʨ��P*��@��B@z(��N	���n��e-����ڋ�"�6�"`�\�;3s��?�o���)�Y��������޽3�Z΅�"0.(Fk G)O�LJ��C���...-..e4��,��J��Q��jW�Uk�T*V*�0���[��r�h�1�6�(b��s㍥r�P,,//��(r	j�^)c֘�GXǎ�c[4H�����(�ƒJ�����Y�-.,�>s��i�*��-���� �� ,��6RHDĝ	�-R.'&&�����̙3�J� ̲�1���]oZ���:I�f�99���}�T)#�4F`�2k���<K3BI�eN��a��� {��u�������Z�Xd�EQ��e"�ܹ��h4�M�Rd���RA(����n�۹\822����G�|��j1�Т�2KSʘ�R�9g��p�HFkJ��RJ�����nm��|��g���iwr�B)������|?�Yʅ���e�㷐�*�p�W���[c�4�����o}l�>cL.�[\\��׾6;; ��SJ��z�V�җ�499����/��"��)�}��=��C��Z�N'�������;�DQ����n�?������KA8�2+�J����⨓��L.�伯\C)�j'��Z�[x�f�LuI!�$���MS�a�1n���k�B�e�(�8KT�ǎ�ib�$iR��a��Z��ѣ���333���O��>24�����������۷��姟~��ѣaz��������������Ϝ�?|�p��i6��68������"�|��׾��3���c۶E�����9Q����"0��[c�8��C
��B@����o8G�p.#�Œ�T��(��������hm�J��Q�9#� �Tie�5F�����Ν3�a�l5WWW<��O�ر��hB��Q'����?��?��W���o���LOO��mkmE��\.玼afY���a����.�������0������>�����v��k�W^y��h4ܖ'�PB� RҞ��J����:u�^�
���99lɳ�i¹������G:��Onn4�����C#�X�*5\0�(���=���xuu�E:666�ǟ���'�4������i��j��k��f�����������nK��R�c666FGG���k��v��Y�ϭ�����w�m���6�Ball�Z��~�\޹s���Z'	%���p���RJp	P'��JQ+�4�͹����P��(�A2���[/�,Zk�D$����ݽg�̍7�Z�0@�QJ�<n,��z�c�W_?|�0" ����f��������0�D���I�8]��ggg�(��ب�j��{����>���=����N'b��cP��lz��|!�ݧ�;44T�V���g���0����Ç���[o�Uk�}�v�4�=�56Ͳ(�.\���G�{�4Mgap��n1���	.�T�Z��P��?�����/~qϞ�CC��\.I�,S�|��;;��#�{��_}5MS�VR�&I>����Z�UN"���,M�<��n9!�@J��t�RRJ�t�j� �1Tp?��Te�Ry����S�Pܽ��8������F��(��F���o~�ܹs��s��f#�������1yuuuyi���?y�G�ΝB�qB���n��b\�"�Et�?��,��J��W_M��>>3s���$�]XX��DQ��Ͻ�����R�fi��b�������ڱCi��*�K/<�⡟��;���;����!�u�ݖR.--���K�ϟ���޺�̌5؉;� o �y���S�߽�n;?;����Z�z���^~y��B.��Q�N�l�Zq�����H)}ϣ�Eq����������o�8�)aY�)e)�ֺ����= ƘV�Ǳ+ʨV�'O�<v�Zmছf�Ձ���z}���\��W��F�4֩�y����b�w:���S�B(�s�	ɤ'e�D�N���ZZZp��R����X�#c2!8m2B9��Պ���fksnv�V-�ٽ������X*�vNNl�>~���o���Ϝ>�$tdd��������V�����\��h4���.�iʹ���qF)G� ��(�Dzi���/��?�����4I)��g�� X\\쇭���'}?���4��V����d���j5�� �IBh�i�y^��i���q!O��k��K�XkA���l�jC�R���m�Z��1�ʥru����Y��gffn���0����V_s!�rZ�ӝ����� �����'���?�#���Q+,!��(s��~��Rjrr҅Ń 0�87�jm]� 8p�ԩ�z�8��h,��J�z�N)�V+.!�p�����E3��0t300 �Eq��i�ZB�$�,UJ���ϟ?/�x���o��j�sc.F i��`bm�����ey��pC�/�y?���,����T����DQ�$�ӗ��"�,K�N�\���7��(��~�qd���s�$�9B֚����� ���2ƌ��\�R�4�M���y��Sƚ�f����o۶M)����$����p��>JV7�����V��x�V�ո��}����f��H ��w��1q��5�U�2.X�B��I[4##��!D�PP��t:a����K!�� ȹpŶ��r�"�����e!$MS)����Z��8��sۄ�I���uDt��.��D�=�7�"}�'�ĉr�\.��<m=^vS���Z�688t~�|���v'T)�K)i��!]Fk!y�X�*�=/��Yc���ʀ�������*MSҝυ�-�$�Z%�gDp^,�6I��q.�`�S���(1��Q\*r�_��:��[��,��3��\���N.�J�R�e��J�����r���@� ���x�>��y'�XHϣ�[Y�0"����BkU� pb|"˲N��$���R�h�q�2D�5c��<�G�K>C�ә��P�T��@�.ލ����ՕV�522�>���n[�ݩ�mg�6��{Z��!c.��4���B��<c��y�� ����j�Ȗt�˳��6NIOh��,}��W�8�|��r��]{�����J�(��B.���0F+�������P�i�0Ƃ���(�1F����T.� Ji���q!e�eBx���SSS�r9�N�s�-�
�����)D��jL?+�g!��}JY��w�q��ݻ��nk�����y;�����?00�^H>��T*n���Ҷ��j�δV�:*��,5Jmj����ʩS����rIJ���������I�y��2I�uǍF}�ðR�������9�J��4BXkj�ھ}�(�+++��������뛛Έ@/z�4��4M�(��J)=)p۶m��w�Ν; I��/w��W�v�~�W������V�������SJ� �<�M�U�J� h|)K�<e$���B�V�n��/���eIZs�2FH����P�I�����y�T����y4&�t8��4�KighC/HӔ1ZD�//;H�����������1���s�P�F��F?A��Y�j�C<����ߟ�睊���r���ww��_���w���s����xE.4�U�$H)�
�s��dY688x�������qI!�$e�j�Y�gf��ڵ{~~�ԩSI�������[o�5�3��?~�R���7�]�v�A
Ƙ���z�Ni�g���8�YVW��)glxx��?��c���3�p)]�g�^��>�O�ڵ릛o���`qqQJ������R�4��1�9s�*JeJ)���̍�R�С�c�Z�L�(N"���mc7ݴ7SI��qԪ�X �nw��>=�cll[�d��b�����</��_�p�R��}�ݜ󹹹'N���,--e&su��y\:�)�}�eB�<�ȣ��ё�U���.�4!fi��;��~�w~gf���^{��}g_z�t��j�`�RkeD�4�㩩)J��y�oٷ}��r�wb��ʨ�U+U�u�R��C�����P�i�T�w����ɉ���;�<���榐�X(�K��驉��N�}�7j���|�R��rܿn���	�S�R�8�����?�裟�^Ⱥ�}]�l��ZBiǜs�I���L2�Xcl�h�d�R`�"�,K�6���F�Ѯ�j��pE�f�s�Ɍ��$�#ƅ3x��N�c�e\X��LJOv:'�J)ʘ�s�������\�^_�=/IR��mL5� �ՌPB,��b�P����e�yzn 鵡]↹O@( �� ���2���. �����>����)!V*�L�ō��k��~.�Tj5k��\[:?�X/���S@����}�Pa����qW��G��I�>��iʽ0nn.,\`��m˗G�mc�"��k��������N�5Z+�dn����";\�<\���BJ'|@�rv�,o *�W�Lz��B0ƥ��s9�4aФV)�2�[CB�T
M��j�F���0̌�����p�m��Y�0�8��ĄKm��!�ފ-�
�؝�H��,,�Lʋ���G.K}��t��+�W�,� �&�{���yK�HX��FIw�-!@�E�(a@(��#�� �s�\pӍ젌]�����R�IȻ���tM��]P�W{	ZG�0�%�x��l��EJ)����Cҵ`G��@]�%v_( ��~I��4G��(��ٵ@��?� �
��`    IEND�B`�PK   'sGTM�2hF       jsons/user_defined.json��_k�0ſ��-M[��ۘ/�csOCF��z�&]�LD��wc�|p0��-���8����N��8#�{-��&�ڀ�8��8��b\奆�o���m�w�Y� =�zcGU�V��3+�J��A^?�}�W�}i���Ҋ�0�uVE�����gI��㣝���N���	�5tvHz��J|��5�:�s�(R�t���e�{��o�$�����<zV;?��h\$�b �q>&����j@<���t�w��(��8
�b�x	�;�7J���іU��I�����Ot�Zs;�`���N/�����q�ˡ�;�X���ꄶp��W��F���PK   'sGT��6  �            ��    cirkitFile.jsonPK   'sGT���.Z  $Z  /           ��B  images/334a8ce1-1ba1-41dd-b982-9eb2c842088e.pngPK   'sGTM�2hF               ���t  jsons/user_defined.jsonPK      �   8v    