PK   7SdT �av�$  �    cirkitFile.json��n$I��_eA�2
nqʈ�[H{�7� 	{�h$�8C��,�X3�h���-�LV1N�c�i�h�4#�Ϗ�FK�=���{>���?==_��<{xz��,��ݟ��~�i�����y�������w���.^���8>_��S��Bلc)E������.����s'Mu��C}>��>�}�����_A�
a/f�Bؗf�B�Wf�B��f�B�7f�Bطf�B���V����V����V�X���,)�Ri��b/�f�Ha/�f�Ha/�f�Ha/�f�Ha/�f�Ha/�f�Ha/�f�Ha/�f�8���N�D���N�D� &���Y�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"zB{�4KD
{�4KD
{�4KD
���kge��f�Ha��f�Ha��f�Ha��f�Ha��f�Ha��f�����,)��,)��,)��,)�EN{���,)��,)��,)��,)��,���v�%"��v�%"��v�%"��v�%"��v�%"���v6��i����i����i����i���^;���^;���^;'_��zy.�_��r�}�rx~x��8�)�x��QNX:a�BDc'l�P:a�¾dcW��C鄥���]����.z6v5;�NX�8�`cװ�C鄥���l�Z6v(��ta�cc�cc��	K����J',]��l�z6v(��t�T <9���'0�>�Ǐv������C`���	̧ϐ��]�'0�>�
�v,��|��.?�m�|���p�`���	̧�J��]�'0�>��v,��|�|:?�}�|����3�?X>��tO ?��|��n8~�7�W��(a�Q�����Ow�����'0��}����O`>ݵ��,��|����?X>��t�?��|��/8~��`����i�C��`���}up�`���	̧;�������O�2�񣟲����G��
�,��|���?X>��t�+?��|��]8~��`�����p�`���	̧���������Owx��a���	̧{��������Ow�����'0������O`>�d Ǐ��Ao���G���,��|�=��?X>����?��|�i�8~��`���^#p�`���	̧]R��5��`����.p�`���	̧�i�������O{�����'0�v����O`>�cǏ�mNo7��G���,��|�;
��?X>����?��|�i�.8~��`���Ncl�Z��|�i�48~��`����np�`������鷯O��Ǘ��9���+¥n��,uq캶�O!����14���2��͗9�cS���;�f��4s��ޝ��?6����[f���m.3��O��6ִ3�������̛���;ޘ{��r��or�T�xc�MNr�o�{����{�;ޘ���r��or�O�xc�M�����2�������^c�MN}�o̿�I+���79�$w�1�&'��7������֙�1�&g^�7��䜉�������;u6���<�������a�;�j=��7���;~9����r-�����PD����ۢ9���9\�C{]q�I×�����o~����>i��[�4|��O���'7���e'i�r�IKk��n�u��7fފ�Lo̽י6ޘ}+�3m�1�V\g�xk�3�ߊ�Lo̿י6ޘ+�3m�1�V\g��1�V\g�x��1�V\g�xc���δ���[q�i����:���o�u���������:���o�u��7�ߊ�L�:�o�u��7�ߊ�Lo���[q���9���]G�M'E�w��p��v��y7�����|<��(w�5�x���;D+Ƕ���jW�:�6���^Z_:a�rҦ��m�r�&_�ؤ��	�4|9_����k���j�4|�X&_��iicM�忘�?7�K�����6���COo����6ޘ�+=m�1�Wz�xk�5����6ޘ+=m�1�F��� �yڟ��<=�}��]0��Иw�)�����BB	�Hg� ����
:�`� ��s�
:=b� ��3.�
:�c� ���B�
:�d� �0�^��Um�lcu[��M)�a1a�[��M)�a�1a�[�N)���@LX��SJa�NV�K��SJa�x7��&�X/�:N)���BLX/�:N)���CLX/�:N)��}�	��%V�)�0<y �q��WX������ĭ�pK)X��:N)����	��V�)�0<�1au���8���m &���X����TĄ����R�^���5qnQ��5V�)�0<�1au���8��'� &���X����$��V���SJaxbb��x��qJ)OBLܷ��כXo�:N)�a/Ą���㔒���:�bu�R��SV�[��/)巙�ؕWzC���*.�a��[�
�ՃU\X��c3\���������ʸ*WVqa���%�{/3�`�8r��Ǟ�L<XŅ5�Q\���W3Vqa��ݛqU0������:�`\=XŅ5�?v{�U��z���>�c|������>�ur]N���w�����B+>����Ol}ܗ����3�>��q`.��C������ǅ�Њ��a����s�Z݋�[7�B+>����'�>�̅V|huo�Ol}\������/||�����^%����2Z��=W>�u�F��+1_V����Ǘ�Њ��󉭏/s�Z���[_�B+>��'�'�>�̅V|huo�Ol}|�����Q����2Z�ս�>���e.��C�{v}L��e.��C�{�}b���\hŇV�P���Ǘ�Њ������ӊN�+����ǗU>�̅V|huo�Ol}|����j�����2Z��^	>���e.��C�=|b���\hŇV{W���Ǘ�Њ���p�m���\hŇV{����Ǘ�Њ��D񉭏/s�Z���[_�B+>�ڣ�'�N;ɜ������Ǘ�>�̅V|h�g�Ol}|����j�#����2Z��N>���e.��C���|b���\hŇV{j�Ķ��e.��C���|b���\hŇV{����Ǘ�Њ��j󉭏/s�Z�9�[_�B+>��;�'�N]>��|����Ǘ5>�̅V|h���Ol}|����jOF����2Z��ޒ>���e.��C�=2]b���2Z��^�>���e.��C�=K}b���\h%�����cs>]�kW�K��Y���umџB����ch��a�TY�M����M6Se��w��B��L��^ٙ*ݭ3U�Qg�,t��TY����uP�2ٻt�k���KG���0�t�i���KǄ��0Y�tg�T��,^:�2W��⥳ se�,^:q1W���ss?u�,^:=0W�J0Y�t�^���K����0Y�tD\���K���0Y�t�Y�4#f�x��\&��N�ʕa�x�L�\��d���Q�2L/�ϔ+;&��.ʕ���s{�\�>��r:��E_�m�O��.͡�n�$�lfM��f�$�l�L��f�$�lfL��f�$�0��Y��T6k^Z�A��d��Z@����ki2Lo���09���&�d��Z@�T��,�^H�a�x{- M����4&����>u�,�^H���Lo���0Y���&�d��Z@����ki2Lo���@3b&����d�,�^H�a�x{- �u0Y���&�d��Z@�d�,�^8��Q����8�n:)�c�+������λ����B�/����ݒJ8g)�]u��R���;tE�c[W�c�����$���KR�̼$���KR�̻$�ʹKRIȺ��ҙ��Y9�T6gZ�A���%�
��)2L�n/(��0����&�����B����
i2Pf����B����
i2L����Ǡ�y�{9�\�>����n���������ˏ����CBa� D�Pf$�B	�a��ABa�I!D�Pfe$�B	�a��ABa�y"D�Pg�L��6W���-Xᦔ�8Yg���-X��h#&�~V�)�0�	��qJ)�֋a��x��qJ)���a������%V�)�0z_�	��%V�)�0�r�	��%V�)�0>��0au���8��G#;���
��R�`���n)��V�)�0>��0au���8�Ƨf&��WX����<Ä����R�4b��:^cu�R
�3P�&�-�cu���8��G�&���X����Ä����R�c����x��qJ)��1LXo�:N)��B���v��z��V�)�0�d��:�`u�R�FzV�[��SJڸc��x���%��&l�&���+PVqa�I�?Z����������
�ՃU\X�~�p�V���*.��w��u�k������y�K\'}֑x��k����u�c���������:�
�ՃU\X�~�\�V���*.�a?i�N��q�`V}&���8.Z��g�}b�亜l����%>�˅V|h�Ys����/Z��g�}b���\hŇV������s�Z���['�B+>���'�>n̅V|huO�Ol}����������2Z��=>>_,��2Z�սJ>���e.��C�{�|b���Wb>����e��/s�Z��[_�B+>����'�>�̅V|huO�Ol}|������J����2Z��=�>���e.��C�{]}b���\hŇV���<����\hŇV����Ǘ�Њ������/s�Z��[���W��e��/�||������|����2Z��>���e.��C��|b���\hŇV{>���Ǘ�Њ�������/s�Z�����Ǘ�Њ��񉭏/s�Z��[_�B+>����'�>�̅V|h�G�Ol�v�9m%��e��/�}|����j� ����2Z���G>���e.��C�=�|b���\hŇV{Q���Ǘ�Њ���r�m���\hŇV{����Ǘ�Њ��8󉭏/s�Z���[_�B+>��s�'�>�̅V|h�w�Ol��|8����e��/k||����j/C����2Z�՞�>���e.��C��%}b���\hŇV{d�Ķ��e.��C��>}b���\hŇV{����Ǘ��J��Y���|��׮��-��ű�ڢ?�PK����,�Ü��Л6Se��l��B�L���ۙ*��3U�[g�,���TY� �����97��e�w���\&��V͕a2x� �\&���	͕a�x�0�\�3Y�tJe���KgA��0Y�t�b���K��~�2Y�tz`�4�`�x�X�\&���˕a�x鈸\&��b˕a�x鸳\hF�d��9`�2L/���+�d�ҙV����⥓�re�,^:�)W2vL/\�+�����z��}���t(�C���ۢ9���9\�C{�^HR�̚$�ͤIR�̙$�͔IR�̘$�̈́IRa�e��%�lּ��������4&���d��^H�arx{- M����4�3Y���&�d��Z@����ki2Lo��}�2Y���&M%�,�^H�a�x{- M����4&����d�,�^H��f�Lo���0Y���&�d��Z@��`�x{- M����4��1Y��p*��.Mѵqp�tR��zW��i�!�w�&>Ie��>��|<��(w�5�J�.���A�m]�ծ*SXT���KR�L�$�ͼKR�L�$���KP�,�I*��3Ie�p�e��L�n/(��0�����&�d���B����
i2Lo/(��@5�����4&���d�,�iA����G>}yz�?��v��������������r�?<ϗ�Ͽ�b�-�
���K[Q��׷x<_~{�K���<�_"d������N`�͔������������������z��/O���Ͽ�����r8�⽩O%k���ț+!v�0L��f�0Lۍf�0L��f�0�#�Y"��Ha��m1R�%�`{�f�0�&#�Y"��Ha��m��-�z���P�F�����Q�F�����R�Fݷ���S�F�����%PO�a\��r�QbB
����v�0.�X9�zZ�Ԯ�e+POK���5��d����%PO�a|6�j%�zZ�ԮƧs���',>PO+���5�������PO�a|�����
��v�0>de� �i�S�F�r ���]#��Y9�5Sb���5PO�a|V������v�0>�g� �i�S�F��.����]#�O,Z9�z� �Ԯ�g&�ķP��P@=m�zj��P+PO���5�������v�"p ����T#��ۤ� �7�f3�	�'0_�O�rzH�X>���~�!��C���	�����?�O`��7��MZ�_�O`�8���7i�n�}Y>���< �ߤ����e���I�tN��'0_�O:�szH�X>���~����C���	̧�)�hځ��B�3�tq��ڇmD�v"0�Є�l+Cڍ��B�s�tiG
M���1�]	L(4�>Mǐv&0�Є�,7Cڝ��B�s�ti�
M����1�]
L(4�>�O/T�>&�P�.�1�}
L(4�c�c�eB����)%�S`B�	u�Cڧ��B�^:��O�	�&�}Fti�
M�{���>&�P�w�1�}
L(4��M�cH��PhB�WG?B��PhB�Hǐ�)0�Є����!�S`B�	u/&C��.��.ڧT�O�h�
M�{`��>&�P���1�}
L(4��=�cH��PhB�7Mǐ�)0�Є�盎!�S`B�	u�:Ú�)0�Є�מ�!�S`B�	�O Cڧ��Bj�:��O�	�&��t�(�VڧԴO�i�
M�}1��>&�P{z�1�}
L(4��#�cH��PhB�Bǐ�)0�Є��aC��PhB�aCǐ�)0�Є���!�S`B�	�wCڧ��Bj�#:��O�	�&ԞMt�]���yڧ4�Oih�
M�����>&�P�|�1�}
L(4��(�cH��PhB�ǰ�}
L(4����cH��PhB�kGǐ�)0�l��xlΧk{�p�ۢ>K]��-�S��}}������ބ��'=3�Oz�f���D�?�e�9~҃4s��wh��I����^���cN@kN�Y�����`�\kN�������\k&N���0�Bk&NO���f��,�\k&NOO��f������4k&NO�0,[3qz�N��5����
X3qz`L��5�G��
X3qz(J��y�h����!��L��ؑ+`�����lk&NO���f���\�Y�f��Ȅ\��L<��˵��.�C�n���o��x���pi�uͯ&�_ɂ��+I�4~%�Ư�@���H�� I���J!J�R���ǜ��\�i�\�i�,\�i�<\�i�L\�i�Zh��5��&`��5��&`��5��&`��5����f��5��&`�X�f�_M�f�_M�f�_M�f�_M�f�_M0�����W�����W�����W����L\�i�L\�if�b��5�z*��.MѵqX�tR��zW��i�!�w��?�#9�ʅ%�p>�R����P}w��Z�m]�ծ*��p���K��aI�W,i�J~%�_I���ٕ0~��%�_�rI�W�\Z�����q��k��5C׬r��5G׬r��5K׬r��5O׬r���RZK�UN�f�UN�f�U����}��y�򴏊��>�~��}���;�1Z��o���M������]���{��N�[E��Y�n��E� :��堭#JQ�RG�:����(uD�#*Q8:�����tD�#*Q�ZG�:�����ZG�:�����uD�#��FG4�/�#���~��K�U�� �0�.e��a�v����_�_������g����'w����ƦiĔF,4�I�{���e��p�|��M#v�_//��/7�.�ֻ×/�l~x�>�<|{�_1�Ѷڗ������/�������O?���/���?�Uo��_/��z�?���O_/�/������Q�Gߢ�o/���q|<����W���r��]������������秿����E�>__�]��o��{��p�r�����?<_�w�_�߉��߯�������ګ�x�;�?����/������:&�&v���������S�/EهOC<�?����U��C�v}�^.e���m��tUq*OǢi���NUӅsd��/���8&����)�f�/�������������������C����:�z��r����w�_���}j������۠���r��l����0se^�_�)o�?�h~P=��ͫ��ؙ+���;Z7����n,G�]����f�̿��ƺ���U�}e�p_U�̴p���W�^ž�o��׏��������'���������~�$���C���sWffn�C��m���
�����2�4�qiz�R;�Wo��i��<���Y��mH���������!~�c�����u��,M{�Zn7��P������H��@��8����f����]���8K2�m)�eh����g��<���Y��m�H��e�s��V:��"��8�4s��nd�v߸�+�H�g���� �:|z�����������o��o��|
�t~j��řC�3;�?u��7]��BB�T����'t?N�.��ݩ�"w�"t��8H�͵*�\�k�}��%���iZ5~F��i�c!�l3W�!w�н��7���o��-���̕y�8?��j׾�D�0�0+�sź�q|�7���oSŲ���+��wF�����❻&�ٶ��ߥ�MB5��ޠ�晦�- ��8KT�o�4���D���fn�%*�wx��D��D���fn�%�yg�kow�\��2�4s��ܝsT����ݨ��R��8O5{�,��B۶�����̕y����҉hۄ�͡�nT3W�fn\���s�J'�������
�ܕy�����Yj?�^P��̕y�����k��)�׷��Q�\����q�j��Y*��6mU��5�0�4�oi��9"i�8[�O��0�i���˪���/�e7,��C��8�����ޕ��z�tou��q~x��eS�Uq�OM�CW���XH���\5�1t?����H���}���\�Aپ-��'�^pO���8��?�;�����ѯ������������7i�k%���k!1K��?ډwH�V*)7�\�W�y3����rVoW�����p+�����-�]�>�J^�t�+�*M/��.��+��Q�U�/0�qu��noW��������a�{�|]묚7�ۅq��������Ux�]���n��:�o�_��'�2�ڂ�Y�䅤k~����'\��_n����,�8��?�/wL�Ӆ�i�p�4�n�&���3��p��W1sm�P����PK   7SdT �av�$  �            ��    cirkitFile.jsonPK      =    %    