PK   <tGTk�ԣ  H    cirkitFile.json�[o#Ir���!�6u���e�l��_�%wk��Z=����wgT�*Y����6��i���c(�SU���������yx�_����W_��t����������OW�oﻧ�������{�����������.�7���WM���?�����]����?������R���|����W��B�,�UH]f�*��3DRׄ�
�k�Q�ԭ�Q��m�Q��m�Q����Q�\��2,�)�R��/�a�L/�a�L/�a�L/�a�L/�a�L/�a�L/�a�L/�a�<���ΰD���ΰD� &���Y�kgX"S�kgX"S�kgX"S�kgX"S�kgX"S�kgX"S�kgX"{�x�Kd�x�Kd�x�Kd
���kg��a�L��a�L��a�L��a�L��a�L��a��5�����������������I�x�l�3,�)�3,�)�3,�)�3,�)�3,��6^;��"^;��"^;��"^;��"^;���D��m�v�%2E�v�%2E�v�%2E�v�%R���ΰD���ΰD���Ή���?����������w��ۧ���?H����A9c錥KY����C錥K]�Ʈbc��K����]���3�.{6v;��X�<�`cײ�C錥���l��l�P:c�R�ac�ac��K��-�-;��X�������ءt���]���v,��|~?#?�]�����g0��C
�v,��|~�+?�i�|��}�p�`�����w���g0��+�v,��|~�7?�y�|����p�`�����w��'�a�����k������3��W3��pЗ8`�Q������g0�� �����`>_���,��|�j��?X>��|�?��|��J)8~��`���5^p�`��������4`�������������3��W����g0��e��G�eE�f���5�?X>��|�(?��|���W8~��`���5�p�`����竍������3���I����g0���f������3��צ����g0��������`>� ��,��|�� ��҃^�����?X>���{?��|�y�8~��`���p�`�����F������3�ϻ���ka������]������3��;�����g0��ԁ����`>���,��|����ڜ^n���-�?X>���w?��|�y�+8~��`���~]p�`���������a�����=�������3�ϻ�����g�n~��p��?u�q�o���U���9�W��X��m~�ͺ9����y��?��+���^����D�lZ8�c�����n��-�p��6���?��,M�h��n��W��`�Mv�*̽�W���7�U�t|0�&;9���ֽ`�M�=*̿�^C���7���m|S��M����ͪ��a�?V�j����޵ͮ=�h��o���_������Zڭ�]�>�"��]����?�i��v�;���Ͽ�EÃ�}>����E��~����_4|��.>_q��M4�yw���`���_6>�{g��fߙo�e��w���h��ߙo�e��w���`����_6>��]�J����7ٹ�t|�7��}�J��o��Z��`�M�3+̿�b���7ٷ�t|t�̿�.W���7�Y�t|0�&�9�N���7�A�t|0�&����Z�`�M��)?���@����<�=<^}��M�|[��W���?W��~!����[�J�"H(�g� �䮞!����(`� ���"H(���J~��!����ta� �4�ǁJ$W�����m�
7���sXV�+ޔRεALX�6��SJi8'1a5ܰ"N)���%Ą��
��RαBL�����cu���8�����V�+��SJi81au���8�����V�+��SJi�� �q���X���p�b�Τp�R�:^cu�RJõ�	��5V�)�4\����:^cu�RJõ4�	��V�)�4\󃘰:�`u�RJõI��;'Ν��x��qJ)�e!&��7X���p�b��x��qJ)׹�K?Xo�:N)��z<Ą����R��������M���X���p�Ą���㔒/�Ƙ�:���8��{1&����:>�T����zo\uXuK����$����W�`5	k�>��U��*XM��}�pU0�
V��f�%��ǮVL�&a�� I\?v�b"�`5	k��H����IXS��/�
�U�j��}업��qU���5u�h�`\�&a�{�5�@�$����{�5��.����.�/�8/	�ih�^sMl5�KBkZ�g^[��К������V��$����5��j����4��C[��К��הhb�qdZ����Ml5�LBkZ_㣹���eZ���Z%Ml5�LBkZ_s���芘蒘ƗU_Vi|���4��N[�/�К����ib��eZ����DMl5�LBkZ_[���ƗIhMC�kD5���2	�ih}��&�_&�5����ܘ��eZ����cMl5�LBkZ_C���ƗIhMC�k�5�ݭ(�]Q��j�/�5�LBkZ_����ƗIhMC�=4���2	�ih�W�&�_&�5��|��V��$�������j|���4�ރC�F��$����^"��j|���4��E[�/�К��{�hb��eZ��z�MlE+�DK�4�����F��$�����A��j|���4���H[�/�К��{8ib��eZ��z/*Ml5�LBkZ�%�m��eZ��zo0Ml5�LBkZ�q���ƗIhMC��4���2	�ih��&�_&�5�����V��C��C��Z�/k5�LBkZ�e���ƗIhMC�=5���2	�ih���&�_&�5��Ȕ�v��eZ��z�OMl5�LBkZ�Y���ƗIhm��&��q�o���U���9�W��X��m~�ͺ9�۹}�Ufz���t�-T���]�2�y�Pe�Wv��Lw�B��~ԅ*3�Ufz>�f��L��m�Z*����֪�2L�m`Z*����6��2L�m�Y*�`&��v�,�a�xn/�R&��v\|��o�����V�z�Y5}:��Ǫ^�S�?�Ի�ٵ����\̚E*�f��ŜI�����ա��d�����xܮn�C�vYog��qY�r1.�T.�e�
���E*?I�T.~��\�-R��e�H��w���������3�e2L�^��,�a2��f��×g4�d�,�<�Y&�`&�/�h��0Y|yF�L����3�e2L���\���d��~ȥ2�T��⹍�Ke�,�ێ�T���MoKe�,��Z�T���\Ke�1��s;���0Y<�h���s�t��&����,�a�xn��R��1Y<�c���,�}���O�����oo����y*��?��w��w����p�!���p�!���p!���p>!���pn!���p�!���p�!���p�	!���p.!���x^�)�\���6V�+ܔRO�1LX�6�xSJi<1�0a�۰N)��)Ä�pÊ8��Ɠ�V�+��SJi<��0q�on���
��RϦ3LX��:N)��<?Ä��
��R�@0LX��:N)���cǱ:^cu�RJ�U��;�J��x��qJ)��&���X���xٌa��x��qJ)��&��7X���x��a��x��qJ)�A&�8wR��V�)�4^�e��:�`u�RJ�Uh�	��V�)�4^g.�`u���8���+�V�[��SJi���a�nr�7�:�bu�RJ�V�[��SJ� c����㔒�?ǘ�:�����R�Z�I�Zu\�����$����)�U��*XM�I�Z����$����U��*XM}�$���qH�&a�� I\'��(XM�(��NZ�!P���5u�>q�*W�IXS7�G��qU���5u��p�*W�IX��`�1�8.	�ih��fMlE�Kd�4��4��4�KBkZ��\[���К�����V��$����{�5�ո0	�ih}�&�'&�5�����V��$����5%��j���4��6F[�+�К����h.,h|���4��VI[�/�К���\ib+�"&�$��e�ƗU_&�5�����V��$�����|��j|���4��&Q[�/�К���Vjb��eZ���QMl5�LBkZ_몉�ƗIhMC�kv57&i|���4���X[�/�К���Pkb��eZ���ZpMlEw+�nW���Z��j�/�К����kb��eZ��z�Ml5�LBkZ��ƗIhMC�=4���2	�ih�w�&�_&�5����Ķ��2	�ih���&�_&�5��D��V��$�����.��j|���4�ޣF[�J2�R2�/k4����2	�ih�g�&�_&�5��>��V��$����N��j|���4�ދJ[�/�К��{jIb�j|���4��L[�/�К��{�ib��eZ��z�6Ml5�LBkZ�9���ƗIhMC��4�u������V��Z�/�К��{jb��eZ��zOFMl5�LBkZ�-���ƗIhMC�=2%�]k|���4���S[�/�К��{�jb��eZ[F��Wt{�����zդ��j���վ:V�j�_k�n��vn�B��޴�*3�dUf�x��t�.T��]�2�ݺPe�u��L�B���ϥY%/��s����0�;��j���s���09<�Mh���s�q��@5���]*Ke�,���T����d��z��o�վ^oVM�����W���7��mv��o�E*�f��ŤY�r1gRki��vuh�<Y�v�;����P�]����r\�\��"��qY�����Gi���O�"���E*?G�T.~,R��]�,��e���f����g4�d��<�Y&�����2&�/�h��@5����3�e2L_��,�a���f���s;5�~�2Y<�r�4�`�xn��R&���-�a�xn��R&�綖-�a�xn�RhF�d��Φ�2L��Z*�d��.�����⹽0Ke�,��q�T2vL�m�X*�>�����/O�����cw{��՗���Ϸ������>�nﻇ�C�x��뷗��_~����'����-��}�W�?~��?t?��O}�}����8�����y{����[ʷ����އ�|���D·)�i8��K��|L�",���9A��D�)�i8��K��|T�",���YA��D·)�i<�-[D�$�'P?(�q�4��r 5Ԁ"�H�I�(PG(�q�4��r �Ԁb�H��(PO+���5�xj8�A�G�	)PO+���5�xv;���
��q�4�_�r ���i\#�g��@=��z�H�5����i�ӸF�rD9�OX|���@=�k��BM���5PO�i�T� �i�ӸF/VE9�z� �4����eQ��6@=�k��]��8gJ�4�i�ӸF�9F9�z� �4��ƫ�Q��6@=�k��k��>PO[���5�x�7�����q�4^{�rW���P@=m�z�H���(PO[���5|�7���5PO���� ����S��u��u�޸P7�g0��|���%�����|�n�^��C���̗�I�.N��g0_�p�&�����3�/�/��M�m�/�g0_���4�
�_��`��MzgqzH�X>��R7���!�c��Kݤ��ď�3���S�'д�	�&�{,��.�!�1ڈ�D`B�	��V:���	�&��r�Ҏ&4���)�cH���hB���!�L`B�	�^n:��;�	�&�����&4��cH���hB���>QM���hB_�@ǐ�)0�ф�!~��dB����)�S`B�	}�Cڧ��F�Z:��O�	�&�uFti�M�k���>&4���w�1�}
Lh4��M�cH���hB_WG�B���hB_Hǐ�)0�ф����!�S`B�	}-&C��.��.ڧԴO�i�M�k`��>&4�����1�}
Lh4��=�cH���hB_7Mǐ�)0�ф�曎!�S`B�	}�:Æ�)0�ф�֞�!�S`B�	�O Cڧ��Fz�:��O�	�&��t�(�Rڧ4�Oih�M�}1��>&4��{z�1�}
Lh4��#�cH���hB�Bǐ�)0�ф��aK���hB�aCǐ�)0�ф���!�S`B�	�wCڧ��Fz�#:��O�	�&��Mt�U���yڧ��Oii�M轲��>&4���|�1�}
Lh4��(�cH���hB��pM���hB�Gǐ�)0�ф�׎�!�S`B�D���c{�����zդ��j���վ:V�j�_e�n��v�ca��Io��񓞂��'�U�Oz����2-?�AZ8~�;�p���g��I����	'`4�۬�
Dsp��Y�@4�[��
D�p�yW�@4��e�
�ka4�;K�
D3q��S�@4��'�	�7�~��T�}�ެ�>V�cU�֩�n�]���s߈�ƟɂE��$���gr`ю�g����g����g�������#�lG���3�E������g
��g���	'`4���	Ds�܌`�@4���	D��܌`�@4���	�ka4���	D3�܌`�@4���	D3q��a�wZ4�{�
�����8�^�T ����J��8�B�T ���M�J��8�&�T <C�f�tG�R�h&N��*�f�t׬�yv4��T�
D3q�3T�@جD3q��R������zx{�������oWKl�՗�W)SX���O�����u���m���1Á~����ǚl~����Ǜ0Q��j�����|D�#*�'�>]-1�S�<pI��?���Q���G�>�p|D�#jQ���G�>����h|D�#�����G4>����h|D�#Z����G�Û����	�-g��1i��'ϙ.�ݣO�_����u������w �����OC��\�Y�]�����>�Uww������ŏ�?��o�C����|��O�/���/���ӏ����?���������~�����M������hW��~�����~��Y���q���O��������]���c��?o��՗�̘c�����q���<���{�����������p��c�;�Se��?n�nr@��m�9Uu�����g�ɶ�!��˱u�?�W�nw\o6����cm�W��Wv��ׇ��z������i�<fIU�t������~$���=?ts�xs�?�:�6����Sմ�>}m��s��l3��^��7��|����j�^�����i�9��޾Z�������p���#��{}���f8��>����0b]�"�6�n^P�4��8�ڎG�^��p親�c/U;�i�/4㑛��?�jV=��_�����������!9}�4���{��8}��_�����O0͖��M���q�|=}ܐ�'��6|����?�~n���1~P�s�lyR�vM��� �n���٥��gǶ��:W��ˇ�z_�����n�V͍mW�uu\��~��ڵm�x���c�[4�YP�V6&�۟\6��]ٶ���CU]�^���3���:�mzY�>�n>[[���o���U���?Dz5M��K~����|���u�W��zw�^m��ꦺ��_��7U�ԹR>�Ӣy�|j�=����D�S������sm��I��u����E�Z�>L�8-��j_��^�O�hv�e��0M8��R���ܼ|�nF���W�5��u�ӯ5=0~��ڝ-˿�EP3����_g�\�,� wid|�-���1�������<���9=p��ā���mZ�-����i��i��q3D��N����-��?t��3/����/l#`�~{���~�wG̼��#N�p����L�-/N<scz�͉OBջ�g�����\�p�v|_����'ߞ?�����D�}��A�__��3��ΰ�8�4T;@�	��t��P�g�Nx������Nc�;b���q�����޼��GN���3����^�}}��� PK   <tGTk�ԣ  H            ��    cirkitFile.jsonPK      =   L    