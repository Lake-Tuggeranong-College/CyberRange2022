PK   �PKT���$  %�    cirkitFile.json��n$I��_eA�2
nqʈ��{�7� 	{�h$�8Cl5Yb�ff��w�[��b���>�
5ИiF��-���{���~�|���qzz���ry����x�Y���?��=���p���q��������>���]����Kq|��ǧ8f_��	�R����E-M]�uS�N���ׇ�|ڇ}���˯�����^�V��/�V����V����V��o�V��o�V��ߙ�
aߙ�
aߛ�
�F��Y"R ��^+�^,���^.���^0���^2���^4���^6���^8���^:�qne��f�Ha��f�HL4���N�D���N�D���N�D���N�D���N�D���N�D���N�D���i����i����i���M����^;���^;���^;���^;���^;���^;�a_�k�Y"R�k�Y"R�k�Y"R�k�Y"R ����Y�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"�{�4KD
{�4KD
{�4KD
{�4KD
{�4KD
�+"{�l��,)��,)��,)��,���v�%"��v�%"��vN$�>���\<�$?���������q�7R���'���t�҅(��N�ءt�҅}�Ʈdc��	K����J',]�l�j6v(��tq�Ʈac��	K?��صl�P:a��~��n����.�;6v;�NX������l�P:a���@xr;�O`>}���.h{�������O�!����O`>}���4X>����]8~��`���'��������O������O`>}���<X>����t8~��`���'��f��|�� 8~��`����p��o8�8`�Q������'0�� ����O`>����,��|�k��?X>��t�?��|��N)8~��`���=^p�`���	̧����4`���	̧���������Ow����'0��e��G?eE?f��
��?X>��t�(?��|���W8~��`���=�p�`���	̧���������O�I����'0���f�W�����O������'0����O`>� ��,��|�� ��Ӄ�����5�?X>���{?��|�i�8~��`��ӎp�`���	̧�F�������O����k`���	̧�]�������O;�����'0��ԁ���O`>���,��|����ۜ�n����?X>���w?��|�i�+8~��`���~]p�`���	̧�������`���ip�`���	̧�����������o_�/�/�cs>]�kW�K��Y���umџB����ch&�e�؛/s�Ǧz��?v���h����;3�l��9�c�����\f�؟27m�ig̻��_�㍙79m+w�1�&'\�7f��T��������;�Z���79�(w�1�&g�7���|�����������e̿�96���������;ޘ��Vr��or�I�xc�MN�o̿�)��3?c�Mμ�o̿�9���79�!w�l̿�y
���79� w��z�o��?w�r�����Z��G�ӡ��5D۷Es<]�s�4����:��/��I×������}���>i��;�4|��On|ߗ�N��媓�6ִ3�݊�Lo̼י6ޘ{+�3m�1�V\g�xc���δ�ֺg̿י6ޘ+�3m�1�V\g�xc���δ.c���δ��^c���δ���[q�i����:���o�u��7�ߊ�Lo���o�u��7�ߊ�Lo̿י6u6�ߊ�Lo̿י6�j=����:Oes�å)�6���N��X���x=��9��np����x8KQ�k|�P}w�V�m]�ծ*u�mxi1��,�t���M{q���M���I×6i�r�&_Kׄ���2i�r�L�\+��ƚv�1In��.-/L/m����6ޘ�+=m�1�Wz�xc֯8����jk,�+=m�1�Vz�xc����A`��?=}yz�����`��1%��K�������
���ABAg	$t��ABA�2$tz�ABAg\$t�ABA�$t��ABa��B%���\���`��R
�b�j�`śR
�\b��`�R
�'���.X����� &���X����� &n��M��:^bu�R
�����:^bu�R
����:^bu�R
�7�V�K��SJax� ��X��:N)��		��[I�R�:^au�R
��!V�+��SJax�b��x��qJ)O�@LX��:N)�� �	��5V�)�0<�1qk�ܢ8V�k��SJaxrb��x��qJ)O�ALX��:N)��I8���7X�����Ą����R�,���o7��7�:�`u�R
�^>�	��V�)%m�1au���8���0&���X_R�o3��+�:�"TŅU\X��c�2\��������.f�*WVqa��ݕqU0����}�K\?�^f"��*.�q�׏=��x��k�����c�f&�����7�`\=XŅ5�?vu�U��z��k������q�`V}&���8.Z��g�}b�亜l����%>�˅V|h�Ys����/Z��g�}b���\hŇV������s�Z���['�B+>���'�>n̅V|huO�Ol}����������2Z��=>>_,��2Z�սJ>���e.��C�{�|b���Wb>����e��/s�Z��[_�B+>����'�>�̅V|huO�Ol}|������J����2Z��=�>���e.��C�{]}b���\hŇV���<����\hŇV����Ǘ�Њ������/s�Z��[���W��e��/�||������|����2Z��>���e.��C��|b���\hŇV{>���Ǘ�Њ�������/s�Z�����Ǘ�Њ��񉭏/s�Z��[_�B+>����'�>�̅V|h�G�Ol�v�9m%��e��/�}|����j� ����2Z���G>���e.��C�=�|b���\hŇV{Q���Ǘ�Њ���r�m���\hŇV{����Ǘ�Њ��8󉭏/s�Z���[_�B+>��s�'�>�̅V|h�w�Ol��|8����e��/k||����j/C����2Z�՞�>���e.��C��%}b���\hŇV{d�Ķ��e.��C��>}b���\hŇV{����Ǘ��J��!���|��׮��-��ű�ڢ?�PK����,�Ü��Л6Se��l��B�L���ۙ*��3U�[g�,���TY� �����97��e�w���\&��V͕a2x� �\&���	͕a�x�0�\�3Y�tJe���KgA��0Y�t�b���K��~�2Y�tz`�4�`�x�X�\&���˕a�x鈸\&��b˕a�x鸳\hF�d��9`�2L/���+�d�ҙV����⥓�re�,^:�)W2vL/\�+�����z��}���t(�C���ۢ9���9\�C{�^HR�̚$�ͤIR�̙$�͔IR�̘$�̈́IRa�e��%�lּ��������4&���d��^H�arx{- M����4�3Y���&�d��Z@����ki2Lo��}�2Y���&M%�,�^H�a�x{- M����4&����d�,�^H��f�Lo���0Y���&�d��Z@��`�x{- M����4��1Y��p*��.Mѵqp�tR��zW��i�!�w����%��_*��-!��%�p>�R����P}w� Ƕ���jW��
I*������yI*������wI*�i����u	*��3Ie�r&�lδ�����K���Sd���^PH�a2x{A!M�����4&���d�����4&���d�,�iA�Ag����rx��}��]7��xM������×󏍇��03@� �0�2"H(3�
��!���0�B� �0��"H(3<�
�l!���0�D� �0�b��Um�lcu[��M)�q��0a�[��M)��F0LX���SJa48V�+�R�Ä����RM!��Ϳ�	8V�K��SJa��V�K��SJat�V�K��SJa| �a��x��qJ)��F0v��V�)�0>��0q+)�R
V�+��SJa|6�a��x��qJ)�O�0LX��:N)��y�	��5V�)�0>i�0au���8��g�&nM�[��x��qJ)��z1LX��:N)��!4�	��5V�)�0>�|������R�c��:�`u�R
�#���&��&V���SJa�E�0au���8����0&���X���qƄ����KJ�M�&M�hձW�*.������*WVqa�Is?Z���������:�
�ՃU\X��r���:Vqa�� ��N��#�`�8Gq���:Vqa�I�uZ���������:�
�ՃU\X�~�X�V���*.��L��1�q\.��C��6����u9�.�%>�K|�������>��q_.��C������ǁ�Њ�>��[�B+>����'�>N̅V|hu/�Ol}ܘ�������82Z�ս1>��qe.��C�{||�X��e.��C�{�|b���\hŇV�\����1���||Y���J_�B+>���'�>�̅V|hu/�Ol}|�����D����2Z�ս�>���e.��C�{D}b���\hŇV�����Ǘ�Њ����y0�Ǘ�Њ��=����/s�Z�C�[_�B+>���'�NO+:=����*_V��2Z�ս�>���e.��C�=|b���\hŇV{%���Ǘ�Њ��|����/s�Z�]�[_�B+>�ڃ�%���/s�Z�%�[_�B+>���'�>�̅V|h���Ol}|����j���:�$s�J���j_V��2Z�՞A>���e.��C���|b���\hŇV{8���Ǘ�Њ���򉭏/s�Z����Ǘ�Њ��󉭏/s�Z�q�[_�B+>�ګ�'�>�̅V|h��Ol}|����j�<��:u�pj����_���2Z��^�>���e.��C�=}b���\hŇV{K���Ǘ�Њ���t�m���\hŇV{}���Ǘ�Њ��,����/s��4�������tm�].u[�g��c׵E
������Y:�9Se�7m��B7�L��>ޙ*��3Uzeg�,t��TY�G����A:Se��sn�A��d�ҡ��2L�.��+�d����2L/�+�d��a��2Pf�x��\&��΂̕a�x���\&���5���e�x���\h*�d�ұz�2L/^�+�d��q�2L/Ė+�d��qg�2Ќ���s�re�,^:m+W���3�r]��K'G��0Y�t>S�d�,^:�(Wf3����r-�����Pԇ:}ݷEs<]�s�4��������5I*�I����3I*�)����1I*�	�����f�KR٬yiY%/���ki2L�n���0���&����Z@����ki2Pf�x{- M����4&����d�,�^H��e�x{- M�J0Y���&�d��Z@����ki2Lo���0Y���&͈�,�^H�a�x{- M����4��d��Z@����ki2��c�x{-�T6G9\��k������8���.�C8�M|����}*��x8KQ�k��B]�ݡ+�ۺ:�]U��$�0,������xI*�y����vI*	Y���Y:�T6+g��f�L�:(y���^PH�a�w{A!M�����4&���d�,�^PH��j0���
i2Lo/(��0Y�ӂ�����-�|����8���sy�ׇ�˷��/���x�?=�/�w���0[0�_��������o�x��������y.6�D�x�?����%����'�)�����ǧ�����%�������:��_����w�����p>>�{S�J֚���7WB�a�v)�a��)�a��)�a�F
�Dl���,�b�0K���)�a�MF
�Dl���,F�f-[D�$�'P?(�v�0:O+PC(�v�0z_+PG(�v�0�o+PK(�v�0�+POK���5¸a� �Ą��%PO�a\D�r ���]#��8V���@=�k���+POK���5��l��J���]#�O�X9�OX|��V@=�k��#+PO+���5�������PO�a|�������v�0>�e� �i�S�F4�rk�Ģ)POk���5�������5PO�a|Z������v�0>/h]��i�S�F�X�r ���]#��LZ9�o�����z� �Ԯ�-�V��6@=�kh�?���-PO��E� �i�өF~�IgANol�f��O`���t�����|���C ��ď��/�'��9=$~,��|�o��^7��,��|q~�o�^����|��y �Iu����	���n�?�O`���tD�����|����9��ď��O�S�'д�	�&�g,��.�!�ڈ�D`B�	��V:���	�&��r�Ҏ&�P�)�cH��PhB}��!�L`B�	�Yn:��;�	�&�����&�P���cH��PhB}��^��}
L(4��]�cH��PhB�wA����ʄ�)%�SJڧ��B�~:��O�	�&Խ:ti�
M�����>&�P�H�1�}
L(4���cH��PhBݛFǐ�)0�Є���~ ��)0�Є�'��!�S`B�	u?#Cڧ��B�^L:���]��]�O�h�R�>&�P���1�}
L(4��ߥcH��PhB�{Lǐ�)0�Є�o��!�S`B�	u�7Cڧ��B�~u8�5�S`B�	u�=Cڧ��Bj� :��O�	�&�ti�
M����;Q�(�O�i�R�>&�P�b�1�}
L(4����cH��PhB�GBǐ�)0�Є�K��!�S`B�	�Æ�)0�Є�Æ�!�S`B�	��Cڧ��Bj� :��O�	�&ԾGti�
M�=�����m�Oih���>&�P{e�1�}
L(4����cH��PhB�QFǐ�)0�Є�_�aK��PhB�Gǐ�)0�Є�׎�!�S`B�"|?d�؜O����R�E}��8v][��j����鉅��'�	3�Oz
f���V�?鉚9~��4s��i��I���񓞟��'�:s�ǜ�����+`����f��,�%�+`����]��L���+`���L��,�+`���YN��L����+`���yE��i�L���+`�X�f��0�\k&N����f����\k&N�h��f��P�\�њ���Cr��8=�#W����32r���L��J�+`���9�f�b���	�+�xn��k��]N�"���o���t������_M��I�W� i�J$�_I���+�4~%��[���B�4~���9���W��9��W��Y��W��y��W�����W�̵К�k~5M���k~5M���k~5M���k~5�3͚�k~5M���l��5��&`��5��&`��5��&`��5��&`��5��&`�!Z3qͯ�	X3qͯ�	X3qͯ�ͳ����W�����W��fŚ�k~�T6G9\��k㰺����8���.�C8��~�Gr2�Kr�|<��(w�5�z�.��͵ۺ:�]U����+)�4~%ÒƯ$X����J��^I�W�+a�J�K�R�Ư���1' �1x�Կ�=k��Y�4k��Y�4k��Y�4k��Y�4s����5��&`��5��&`��W�����������i��}��.e���/wZc�.���*�[���o�����o��7Ꝣ���+z��ݢ���/:@tD�#�A[G�:����(uD�#JQ�JGT:�ptD�#*Q�JGT:�����uD�#��7����uD�#jQ�FG4:����h�_ZG4:����z�2����	`�]��=vÀ��!ؿƿ������E���+��O���O�Mӈ)�Xh���"�r������x����F��_^�I_n�?\�w�/_�?���x}�y����b�c�m�/�����e_H�����՟~$�G_.��Ϋ�"��/��z�?���O_/�/������Q�Gߢ�o/���q|<����W���r��]������������秿����E�>__�]��o��{��p�r������?<_�w�_�߉��߯�������ګ�x�;�=���^��_��uL�M�T��ӷ�����_����x�}>�8�V��5���U{���#�?����Uũ<�����:UMΑ)~��O㘤������=�F���_�Nϧ/�׷���^�����?�ݧ^��_i+�Vu�O��_�p�4sa^`W���x[_�f��K4�K5�����G��yU;s%U�|}G�f���ˑf׿�bw{��+�5���?��G�x_�,�W�?3��-��nx���w����w�����������'���������~�%$���D���sWffn�e��o����
�����2�4�q�iz�S;�Wo���i��<���y��}L�������)~�c���a�u�N�Y����F��PJ;�P��Aw�z��<���<���P9"w�(n@sW�	�7ΣL�[`
s�����=��2�4�q�iz�<��|�o�ѹ+�L37�2�ܷ������n��<���y��}3L�������^�������m���O��U�3�8�h�qfj��.V��k^#^H��vW�����)�%����J��S�K_�n��Z��J.ݵ�>Nْ,}Ҕ�?-o����8'��R�S��5e�1~��}��oy_�$f��KĹb�W��uV"7��Y�7�}��k=�	�\�x�6�͇8�]I��v�3Z�ח���5�ζm��.�&���oP��L���fn�%��7d��y��}D37���;��G��y��}D37��4����I.�\�g��qj��9�a.�v��nTsWf��n����s�Jg�m�To
͍j��<�̍Tsw�R�|�mB�fVv7��+�T37.P��9K���x���sDn�v��<�̍Tsw�R�L���a�	(Սj��<�̍Tsw�R�5~���[�ݨf��S�ܸ@5w�,�N[���߂z��^�g�޷�4s���e���'�x_Ҵ�T�eU�덥�Qv�"�?�����ٽ��A-^���wM�V�����\6U_����1tũ���T;��UsC���0�k����~��ǉk̕���۲�.~���Ԩ���c��S��0�M1ʺ���R�Oޡ��k��8���V-@{���x��㡝x��o��rC��}�7�����+g�vEK�^i~X�
�R�?���*�ەq����uLw�2����Z�By�2."u]���ZWw{��ve\���h߯��V�w��eϪy�]�r������\�7�ۅq�_�v��Zw���~2,��-x�5M^H���/]�y�~����	���.�����p��=]�q�7N3k��ir��8��73׶
��_PK   �PKT���$  %�            ��    cirkitFile.jsonPK      =   �$    