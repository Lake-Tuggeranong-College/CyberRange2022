PK   �\IT��v˘  ��    cirkitFile.json�]ێɑ���u52�R���1���mx�Q$�3Ķ�Z6{f��|�f�i3�lu�2�*�qJv$��R3�TDƩ�fU��8�?t�����-���������a�c���f�aw�<����/���]���+�������qiպ�ݦ.Vۦ)l�]mY�4u�蒶۪\�ś��n�6'��������;�y)3�d�̼�&�.e�YmWMٺ�+�+l�^+S��z�Zw�δnC���KS��kM+[wE��v�]�MQo[��UUn�Ҷ��K�K����C��[��N���­����m�ƭU���ҕi�̒�������;�����"�wHx���!��C����7	� -��t��Z�?-��O����+�ږ�F����]��vd��6��̚j;2o����g���2��e�O=�<�y�y>�,sa����<?��h#���w$$�ȬǳRod����72������x㎐#��^ȿ�Y�g/��Ȭǳ�O:�i!���F�?#䟑N�B�!���F�?#����g���B�Y!��t�'���
�g���B�Y!���N�?'���I�B�9!�\��*��_Y��x{��Ӷ�t�荪Und��2�g�e�O>�<�{�y>�,�|�Y��ĳ̅y�;,���ã��vBލ�:y�B��:y�B��:y�B���:y�B���:y��qOȿ�]'�^ȿ�]'�^ȿ�]'�^ȿ�]'o��od�ɳ�N�B���:y�B���:y�B���:y�B���:y�B���:y�ҕ��#�N���#�N���#�N��Yȿ�]'�^ȿ�]'�^���odש�vk�V��{M��,ںm�v�l��f]�����=�s��J����I��G��̶j6Ū"��.�m�j�*�uS5��6몕w��t��	����q��L�W���=3��4︒�����16}i���ʫC�nV����1VEb�k9��)�a���w�%�k�#q|�����H�{}�6�͟4>��G��T$����56�?i|�����H�~}�l�6��a�S���p�͟��Oa�#l|*������s��I�#l|��OE_����Kl�Jl���6>�Ƨ��,_��66��a�SїƯ�����?i|������[��wx��_�͟4>��G��T|l�7X�!�#��!8D^����:Z�(1h)&
�zWu����+9�r�!8D���C`W�:X�!��#��!8DŻ�����eq���!��@���v,�C$p�Q��R��u��C`�G"�C$p�*>|E��u=�	"�CT��+z��X��H�	���_��`͇���8D�H�U����ԃu���5�W�r�b|>Op�M	��y�+��4X2�H�	��������x�'x Gx�gx��O�����}4X��H�	�����������>�	"�CT�s�W�:X��`�G"�C$p�*~�^�>,��C$p�Q���^��`�g���8�r�b�$����&E�i�b����8D�H�U�h��V�4X1�H�)�/=`x%�z�?_	�����,n�F!������8J	A� (5����'����SZsb���#	̙�����/aL��0aHLk��Ac0f�k�5���b=�b�K�(���"�2���(���>������}�<�u �b�K�N�����#`0�����G�`H<=s�_P����O����#`0,����o�G�`X�1,6�h)�a����`Xl0,6����b�a�Ű؂V�[�-���b�a�Ű�aX�0,v;�hc�a�ð�M����~ �$k�/��Lr�� �$c�/��`�29�q��`���Nk�* ��� vi ���Z �^ b�ðxZ`@�`X<��+ `0,����0Ok��R��i-�]� �a��.Z����xZ`W2@�`X<��� `0,���50Ok�B��� vuhc�a����P�燸E<
)UVin�q_���i�U��6�­# @�<��}����3��S9���)��_�G�O��P�z?½���pTX�*���_�Gft��~8*0ә�V�B8*0Ӡ����Q��ά�����3
:� Gf:�\�	��3
:� Gf:������3
:�1 Gf:����3
:�F Gf:�.�K�Q���-��3� ����L���+�Q���h��pT`�AAǵ�H�&�E��H����w�x(�8�l&�l&����$���~�p]�Pb�Q̢��|�4�Y�NU ��0�,�?��E����w��(�0�,�T��E����w�P(�0	-�i��E����w��(�0!-�~��E����w��(�09-����E����w�L(�0Q-����E����w��(�0i-����E����w���
L_��4�a�GV`��,q'�T`���#J��xXd�a��,q'jR��o܁��N��t$w&m�Ci��k��� �,��|���Y�NԹ ���E%!��|���Y�NT� ���E�#��|���Y�N�� ���Ee&��|���Y�NT� ���E)��|���Y�N�� ��`�ZT��7L_�%�D����עJxXd�a��,q'
u|�}���pl���^�}�x<�w/�}%
AP4�@P,�APJJA�!(�u �b�K����!0aL
�Ä!1aX�1,֠1�b�a�ưXcX�1,֓,f�됣L��]�C�2�v�9�$c��:�(�Lz�z ցȋa���ͯ���xz���� �`8<=s��u F=��gn~� ���37�^ �b�̭1,���������`Xl0,6����b�a�Ű�bXlA+b�-���b�a�Ű�bX�0,v;�����ð�aX�&Y̮�!G�d�^�e�3�zr�Iư�u�Q0|����: ����i-�_� �!������pxZ��� �zOk�z ��� ~� ���Z �^ ��i-�_� ZJ`X<���u `0,����: 0Ok�z ��� ~� ���Z �^ ��i-�_� �a�����m�0,����:�(��f�됣L�®�!G���[�C����z	 @�4�� + �l �:Ш��U�2�zhT`�AA'�u�Q���L��zhT`�AA'�u�Q��ά� �:Ш�L��N��@�3�Y��u�Q����ׁFf:�� ��@�3
:Q��
�tf��ׁFft�^�錺�ׁFft�^�� �ׁFft�^��F�ׁFft�^���D��n)��t�Y�N����'�ͤ��$��Բ��y��܉-D�8,2�0�l��S�:0���fq�
8,2�0�l��S�:0���gq�
8,2�0�l��S�:0��Ihq�
8,2�0m��S�:0��	iq�
8,2�0-m��S�:0���iq�
8,2�0Em��S�:0���jq�
8,2�0]m��S�:0��Ikq�
8,2�0um��S�:0�U`�Z\��<���f�;U��o��׭��"���f�;U��o܁��N��t$w&m�Ci��k����:��|���Y�N�������u+��|���Y�N�������u+��|���Y�N�������u+��|���Y�N�������u+��|���Y�N�������u+��|���Y�N�������u+��|���Y�N��x��������r������O�7�f����=,?ܵ�n���/��MwX�y��ى��J�M����-V��¶��MGMQ�n��%QK�e���V�sm�
���®�T�[S�Ѷ�kgJ�Ml��ݼE��\]��l���7ОN+ohU犺6e���r�ve����W�c,�^�ᒽ+�+��ēWf>�,������ǫs��Ε\>xO�g��|2>yen�ܥy��.=��Ō�M����f����ƙ('���ݹ�q�Y�2��%MWn����v(�
���d�wO��C�~��_����J���7����ϯ?��������~&<�̻�ޣ/���Y��#�ɣ_��/G� �7`�"����Ac�3�y<����B�;�V�F=�,��#�N4��'���=��Q/@<�H_�Kc��繣�Zk��S�܆i�C���1�}����r?E�$�?��:2T}:�	��s�[p\��z���]���'�qw�_>�c�x������t��q�|�mo~������R�V�k���[��ڗB�Jh_�)��'[=GxV��c�R�'%,IKRʒ��$%-IYKR�j鸩��t��R&j)���Z�D=�DVm���GH��,,�� ����~� ,{i�G"���8�㏘�R���c3"@J±� ��،��qlF�DR&�͈< )�fD���c3"@�D񌨥L�R&)���F<-K�h�L4R&)���F�D#e��2�J�h�L�����V�D+e��2�J�h�LtR&:)���N�D'ެH��Lt#Ld�a����~���B�
��X
�G����d bُ�C<��	(e��~� ���~� e��~� ���~� e��~� �Lۯ� �Lۯ� �Lۯ� �Lۯ��4)���< �,e��~� e��~� e��~� e��~� e��~� ^!J�8�_�H�8�_�H�8�_孳�Lۯ� �Lۯ� ě)���̳c����h���.sΙy�,����w&�<��㟋a�/��a>1��׿(@^�����8�ӻo��I"�C$p�*֛�x�98����Y�H�	��U�+^��b�^`a�!8D��b�������ɢ8D�H�U����ףW��� Y�H�	����x}�G/���A�(��!8D��^�^��ÃdQ"�C$p�*�N����L�ɢ8�D�{$�����^�^��ÃdQb�|=��Hw|}�G/���A�(1Q�����ě� ;���7�(S祹DH8p.� T��E9� �U奙@;qEuij�8�T�x�m
Pw��@@L.8�TMxi.O\��%@�G���.�%@�k�1��=�(S�ܥ��=qs  &� �e�N�4� �'�Q�� ���L�`������ǁ��\�p�����\���8�K��2U;]zl  �uÁ��� e�.��A�+�K3�V������T!p�����q�~�~�q�~�-ŏ]��h(.�-�%@G�*].�%@��v1��@�(Seɥ��@qIn  &� e��4� (.��� ��L��� ť����\d p��R�-
	SP���@@Lj�8�TUp�m
P���@@L.�8�T��e����|�n^c���c�ym����Ex:,��A��Ņg��h�HC��_��7�M�0����N�-��ZShN�=
:X�;X�`���:X����=_���?�B,L�0�;��,L�0��,l�����G,l����,l�p����؊�:X�`���<����.�6���s�y�#���J/z�0�����޿���_�=L���W�=~ 7��'�^?��v��4����x�Ij��k?k��c�\@#xM��T`ڻ�S	�y�8v?�w��E<L,���	�ߴ�G&�Ȟ?��G����?��G�������Q�?�����ow��/�v�����G�Y������a�w��&DN���޺��XZr��牑�}��{���&���_��������_��p~^��|8v���}�>�;|z����{�2��������{�~��_���Ao���C�?|���=�Vw�����y������;�����ܶ���!S�_�e�g7~�i�����?�o�M� �ʻ�W��n�;�mA�{��t�<wrsӸ��ou���������<��5Ͷܮ��8r���!��Q����W��Y���������~}�a��o{���=y�x�����w�9����r����w7o]�Z��Z�o���4��o�=���LCwB4���Z������	�v�vuշ#s�r�¤z��>7��\C��X�:���ο̺H�G4UsF��X���=�N�]u�O�͵kNx�N�6:�g�������=�vY$sB��(�0��\6��t����]�n�,�.&A�]̪d����f1��7Q�]�L�K���h�q#n��n�{w����f��Gwx8�Dt�n�O��iE7�6�W2����u|=�'Ucʮ���U�*���M��땟T�:�����f8����|r��_��n
=�._-��N=�Ͼh�s�:�4��i����ҋI��p��>_�f�Rӈ�AP��3��d�ν:U՜�0��$�/�hHZ��0zT�R��{'�F��m�l���c�Ű�G��s�����^'Z�>M1����m�aګDá[�&�NS�q����h��+�p�W�����J��8�e�J4L��h8�+��үӔM�$�siL�Kz�h7p*�b��	�9w���H��n?��~g��t^�5e�K풾'�|O���ݝ����C&ס��I�Rn%�\�eO+Zu��2w[$�%�J�8�jq�>/��wME��;�0=�%�J6ܫ'�My�r�s�j�a�^M4ޫ�&/��}��w��/�k?���4+��!�5�ۛ��NSY�K*ԪZ�%�
�5�5���&0X_5��eb��T���Ge�����[��-r�U�v��8�ѥ�	㭩J_9�ѥ��������8�ѥ����iQ��ʩ�&�Mݷ0�q�&V�۰�,������~K�'ɏ.<I�x�j��:u�S�ѳ#�O.��݈[d�(��U���H|r�E�`�E�"�EX�����"/�\z7z��x�e]����~�:����ҏD��#�&O�ҳ,���by�$�ѥ'�COM2���f�Ty�"�}�$�ѥ'�COMҞ��oX5QrR�\��h0p#�"�EX+�~�x��sw�>��"�`�E�Eڋ�4�#��`�<�%?��#�b�H�Iړ�_�<ms�s�$?��$�b�I�I�}K~گ�dŒªͧU[m4}��ֿ���կ�/A���a�n|8�5���[*�*l���R��/��K�Zo��hCźrۢ#��V��b�U]M����.�X'RK,$,� ���z�V��_)��ǟ�#~������#O��Ȳ]U�_v�b�\[�<�u�tE�u��E۪��u�A
k��T�gv\G��u���/R��?������>&D+�1���A.B7����m�����ߪ?FV�:��UMC�����w�a�wx����ٟ�V��p���!��C��V���~������N�T�_�'h��Ϗ�W�᛿l��}{�y�o����N�wS��?�lݏf��I+�2?y���P��
�Vƶ��պ^�vHR�	�!I��?�<=�X6�����������W��~V��k/�!�/�@搿�D��=y8�(=��7E�&����PK   �\IT��v˘  ��            ��    cirkitFile.jsonPK      =   �    