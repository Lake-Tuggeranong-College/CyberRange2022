PK   ^IT�<w�&  ��    cirkitFile.json�o��8rƿJ�mX)��.Hp��I$�7�� K�]#���g����aI=ݶ�?��S�n��ݶY�.�K*R,~?\ڟ��{����������#��������������񹹾4��_�r����;���ː�.C۟^�MC�ɇ����8�3K�͎��g�8�E�z���4�����߮@bӐ�A�`�\� U0M!f�*�Ɗ�
�qb��iJ1�T�4��A�`�Z� U0�Q� U�9J�(���*幒��R,�)��R,�)�	S,�)�)S,�)�IS,�)�iS,�)�S,�)�S,���S,�)�S,�) 7��ܙ�s�X�S�s�X�S�s�X�S�s�X�S�s�X�S�s�X�S�s�X�ׄ��)����)����)���2]�;y�Kx
y�Kx
y�Kx
y�Kx
y�Kx
y�K���s�X�S�s�X�S�s�X�S�s�X�S &9���s�X�S�s�X�S�s�X�S�s�X�S�s�X�4N�;��B�;��B�;��B�;��B�;���D$ϝN�;��B�;��B�;��B�;��)�S,�)�S,�)�3�����p�.��S�S͗����x��7����ź����<���t��ʝ��$�ٚ\��C�]�S]�|�y���<�y�|�L^��Y�Δ��|̎=uYo:s�������"
���>��O�E����!?�&�p{����C�JGX:�X�X�A�K���,�wP:�������wP:������J��t��3M��]�����t�����������4G��X�A�K��1b�GQ�L\i%-h���>��W�[�{=He�.M��	��W'X>���`��+,���Y_���U
���|��2��J�G`>~��?p���#0?��b�����i�\�`���O���\�|��}��i��=����; ���X>�����Ы#��p����\`����e���X>��N�������|�G	�?p���#0��\`��������X>��6�������|���������w���?�|����`���,��x�&��'�Џh��\���G`>�-������������?�|���`���,��xo5����G`>����������c�g�����|��?p���#0� �\`�������X>�q���лD��D����\`��ǽ2���X>�q��������|ܟ�?p���#0wV�\`���=a��s���G`>�f������������?�|��B`���,��������G`>���z�:z�:��p��Á�,���S����G`>��������������?�|��jX�����G`>��������{ف��?�|����ݡl�U����2�W��t쩫�%��,�c����-��}S��O��J��-F��A��M=���8S�Fv¸�9K�F^p�X��0���R�����j/���ܪT{i��_p�S��0����R���f�j/������0��S{R�^a�gܤ��/8W&�^�Y.�����OI��_pfI����O�	����N�H��_p�Eꭳ0���#R���ؐj/-=���o�j/���L�T�����i��dո���Q��qe��Q��Qe��Q��1e��Q��e.؍�9�^wc�,�T�7픰�x,�%�e6�,A�$6��8{�b�����,6��8{i:��:>�^��7��8{a�m���ڡ�>�Ҵ��sVS7dy}�W��v���u����e���G���Q��_}���7e���G�����e��u��Fv¸ۘ���F���u��0�6�zq���۸����o�g/�{��۸����o�g/�?�Uoc�:�^��q���ۘ�������u��0�6f����1{g/�����8{a�m�^��K����1{g/�����8{a�m�^��:�oc�:�^��q���C�ב���p�f#ϼ΢��<E�R
���~Q��Kӽ<�\����O뿡�?����o"���oC2�b�@B�'40D !�s$"���iH��L�$dxrC2<߄!	������8+J����K۰�M�čR2� �	��	��QJf��1��7�8JɌ3� &X'XG)�q&���9,����8cb���n�ay<��q��g�AL�<���8JɌ�
 &X�ay�d��,��<�R2�*������QJf\M1�fRpS)�<^��8JɌ+i &X/`y�d�?,��<�R2��$�	��-,���̸�
b��q��(%3��ps�IqX��<�R2�*7�	��-,���̸b��q��(%3>5 Z���q��(%3>� b��q��(%3>�b­n�7ay���8JɌ�'AL�<�`y�d�}� &X/ay��-�`L�<^�����x�W����c?.f��L�X��EV���0~����x d��:�W�U��TXM3�hW�U��TX}ݥ��y�k�4XI�����u��VRa��(*~����x@��TXM3�W�U��TXM3�W�U��TXM3�W�U��TX﻾ ;o&��Thi���B�^Yu)�]:u�^�Sy�В-?k��[��K��th��y��T`*��C�����V�
S�%Z�à�[�JL��thy/��ou�1Zҡ�=%:�թ�ThI������V�*S�%Z�㣳��Q�-���^%���e*��C�{�t|��"��$�S��:uY�S��В-���N]�BK:���OǷ:u�
-���D���e*��C�{+u|�S��В-���N]�BK:���UǷ:u�
-���]��t�2Zҡ��:�թ�ThI���P��V�.S�%Z���[���Wԩ�
���Щ�ThI������V�.S�%Z�1��[��L��th�W��ou�2Zҡ�:�թ�ThI��{W��V�.S�%Z����[�S��В-���N]�BK:��EǷ:u�
-��ro���e*��C�=jt|���Li+�N]fu�2�S��В-���N]�BK:���HǷ:u�
-��r'���e*��C˽�t|�S��В-��R�ө�ThI��{���V�.S�%Z�q��[��L��th�W��ou�2Zҡ�s:�թ�ThI��{���V�ˇR������eN�.S�%Z�e��[��L��th�'��ou�2Zҡ�ޒ:�թ�ThI��{d���ԩ�ThI��{}��V�.S�%Z�Y��[��L���hߏ�n��CUg碣���);��.#{�sI�)��s�UVz�&��t�MTY�㝨��y;Qe�Wv��Jw�D��~ԉ*+�UVz>�F(x1ѻv�k�&~׎VM��D����2�^;&4U�k�q�ʀr0&��N�L��D��Y��2�(^;q1U�k��^u1Q�vz`��V�k���`�x��TL��*��ⵃ�Re0Q�v�Y���k瀥�`�x�TL��i�Zu`�x��TL��ϔ**�0Q�vpQ�&�׎J�ٍb�Y�+w���LfkrY�uv:������P��L�1e%Pٍ�(���Rٍ�(�� �Rٍ�(����Rٍ�(����R�����D�&z�L�q��`�w���!J��D���D�&��g&�d0Q�?3'���$�?3'�I��3q2�(ޟ� �E�����lם���!��S_�µ�k���Tv�&Je7h�Tvc&Je7d�Tv#&Je7`�T0���Tvs^\ԁ���k
q2���_S���D���;N��W�8L�_��d@9��W�8L�_��d0Q�r�)��`�xM!N��k
q2�(�_S���D���B�&����d0Q���'����5�8�1&����d0Q���'����5�����k
q2�(�_S��v�(�_S8�*�W�sV�3ev8�cO]֛�k���=�O�G���\_����寣Ls}i�^��p���]6�{3~������>��
JȌ�����}HȌ�1"���v D !3NA�@Bf�r����8}!	�q*B2��$d�):L��em\چ�m�%n���f"1L��M��R2�)�	��	��QJf���0�r8��8J�L��&X�ay�d�o��w��9,����4��a�����QJfZr�0��x��(%3-�`�`y<��q����i0�8,��<�R2��	7���J�����QJfZ'�0��x��(%3��a�`y���q����1L�<nay�d�UO,�[XG)�i=Ä��M����q�����1L�<nay�d�q,�[XG)�i�������QJfz� �����QJfz�Ä[��-o���q���v�b�`y���8J�L{V1L�<^��8J�����`y����5���rA�B�����J*���j��i!Z�WVRa5Mа�
��+���&h"�V�U��TX}ݥ�נ<������T��x@��TX�=��_���h��
�i���hU�_5XI��4A�x�*Я���j��Y<Z�WVRa�g�u
��K��th��f�*U]Je�N�E:��T^*��C�Ϛ��V��R�%Z~f^Ƿ:�
-����:�թ�ThI���0��V�S�%Zދ��[�jL��thyO��ou*2Zҡ�1:�թ�ThI�����,,��e*��C�{�t|�S��В-���Ҋ�Ғ�N]���e�N]�BK:��NǷ:u�
-���^>���e*��C�{u|�S��В-���N]�BK:��GTǷ:u�
-���^W���e*��C�{vuLҩ�ThI�����V�.S�%Z�C��[��L��thy/��o��VTz\Q�.+t�B�.S�%Zޛ��[��L��th�ǀ�ou�2Zҡ�^	:�թ�ThI��{>��V�.S�%Z�]��[��L��th���o�N]�BK:��KDǷ:u�
-��rO���e*��C˽]t|�S��В-�����N2��d:u�թˬN]�BK:��3HǷ:u�
-��r�#���e*��C�=�t|�S��В-����N]�BK:��SKŷN�.S�%Z���[��L��th�Ǚ�ou�2Zҡ�^m:�թ�ThI��{���V�.S�%Z�[�.Jm>t�2�S�9��L��th����ou�2Zҡ垌:�թ�ThI��{K��V�.S�%Z��R�.S�%Z����[��L��th�g��ou�2Z��}?*�l�U����2�W��t쩫�%��,��aNTY�M����M6Qe��w��J��D��^ى*+ݭUV�Q'��t�NTY���u���D�ڡ��2��];Z5U�k���`bx��TL�ƙ*���(^;�2U�kgA��`�x���TL��k�z��D��適2�[	L���*�����Re0Q�vD\�&��bK��D��qg�2�;bL���*���ӶRe0Q�v�UjՁ�ⵓ�Re0Q�v>S����D���E�2�(^;(Uf7�Mg���)�K2���em?���躞���C�?3���Q*�!���Q*����Q*�����Q*���������8L���L��`�wf"N��3q2�ޟ����D���D�(c�xf"N��3q2�(ޟ� �E�����lם���!��S_�µ�k���Q*�Q��4Q*�1��2Q*���0Q*�x�MzQ*�9/.�@�����+w�&~���q2�޿r��`bx��'����+w�(c�x��'����+w�&�AW��5�8L�)��`�xM!N��k
q2�(�_S���D���B�&����d0Q���'�#�D���B�&����d0Q���Wu`�xM!N��k
q2����k
�Se��t�
w���cv��zәcm]����">Je��R���}����צ{yz�4��_�����e��|yj��o���K?\?}z���-gO/�teuκ�Tg����t�{����b����y/|~@����0���ۇ��1�ܡ"�\�2?�q�%2<Q^����)Q�Od����}���'}~z������~����3�n~�f�eq
�//�$3=$�=��?�e��s"��7��RN�r i���^�o��/��k{�-ӏ�~9�'����|{������2���ŏ��6�ts��*Ar	3�Y
)�f�3R�%̸<%�K�qyKH!�0��B,a��5!�X�sB
�����b	3.
)�fZ^��-D�D�O@�$@�k�i�T�ȡH�r3��J9 y� �T�a�Ub) � ��5̴N-� ���O�fZ)�r �G7��|��\�L��R@>��T�a����|��\�L<H9 �4�S��������|Z �\�L}H9>�����O�fznE�ȧ ��5��䌔�O@>�k���) �Z@>�k���!) �Z@>�k���%)b�1i
ȧ�O�fzK�ȧ�O�fzL�ȧ�O�fzM:�ȧ�O�fzN�ȧ�O�fzOʁX�B,C��S���:H9 ���\�L=��|Z�\���8 ����PC�T�ǃ�������E����	�<�%�n��v���< �B\�ĝA�[��X>�&8i�����|�8�/8FD�y�|��7#`�G�?/���|����8������4��8=���|�3Mp�N�?,��L���Ӄ��G`���w 7� ``Z �z {�/�)J�U	�,!t]B��LHhB~.�Ctq&$4!?Ӌ�!�@���GF�]��		M��R�}�.T���&����>D+`BB�3�h�0!�	��{��E��Є�w =o��MHhB����!�N���l�}_@�����]���:LHhB�+��!�N�����}��S���&�=Jh��0!�	yڇ�:LHhB���!�N�����}��S���&�=y��C�u
��Є���Ct�&$4!�D�]��		M��8�>�?��]��:�@�)`BB��Y��u
��Є���Ct�&$4!�[F�]��		M�{��>D�)`BB�~q��u
��Є���C��S���&�}�h��0!�	�� ڇ�:LHhB�!�N��{;�}ߘߙ��S,�N��:LHhB�!�N�����}��S���&�^&h��0!�	�ڇ�:LHhB�!��C�)`BBr���u
��Єܻ�Ct�&$4!�B�]��		M�=��>D�)`BBr�'������u�C�)]��		M�}��>D�)`BBr�0��u
��Є���Ct�&$4!�f��D�)`BBr_9��u
��Є��Ct�&�=�����v�P�ٹ�(�}u�N��Ȟ��\Ro�"<�0�>�k�h�#L���&��T�>���A��D���h�}�/4�>��?� �F`xD[��4�C�R�QC�* ����Ti$�Gm�
�s�4�S�R����* ����Ti$�g�^Ӥ��.�* �,K#1<�'U@���7��H�I�Fbx�K��4�UR�w��H�I�Fbx�G��4��5Rﳥ��h�* ����Tq�"���Ti$��
lD��,��;e}I&�5������.m>�c�<k�hrae��Q�Ae��Q�!e��Q�e��Q��p�*���8�[MPS��!9��[�R��Ict����F�Vy' �ӭ�:N@�)��r����&˭�:N@�[�5�v(��Ϩ4mf����Y^�����]�5�e�Q�Ae�Q�!e�Q�e/��7Q��F��q J#pk�9N@�[�q�(ܺ"�	H�p�' �ĭ+b��8J#q�' �ĭ+b��4�Wĭ	�8i$nM8�	H#qk�9N@�[�q�Hܚp��F�քs��4�&�����5�' �C�F�քs��4�&�����5�w�-�ĭ	�8i$nM8�	��i$nM8�O�ɫ�9+ܙ2;��ٱ�.�Mg��u}�fk��(�+r3g��ׇû�c�\_������!f����Ӂg�x
��Je>����[�+�o��=�q �$J<�x0�h�����-r��Gm���"g��-r���"g��-
�(آqآ`��-
�(آ`��-,[X��la�O��-,[X��la�±�c��-����±�c��x��p����=��3+��R~���o��.�gx�����m��=W��5~ G�|Fٛ	��o�F�c����C:щ�X�H���Ȭ���2\!����Y	�d���2��_��S{���2�>\���-��%
_�__�×�ח��%�����f���ܜ���|~i��^�eQ�秷���|����۸�)���|�o���-޾����^9������/���8�w?}y���/�{������g���'�o~���s����0cn����Q��}���/����^����>}��_�˟�>�����]����x��ǫg�>��}�vn���p�z��a��ҷ�˷��?����6��ȩ<���<^_�C>eT������9;�.f�?z��)NC�Y[YU�efε�ʪ�S������o���s7�D݈=^�|����������=��ꧬ�?���3�>eu���b�?^ �߿b�^��ݞ
/6�����{;�|U��ި�^��I��>�vo��+gm������z�̋War�_��+.��S�x��yY�x�)	��P��M=���.?���(^���:_�H��>`为
"py\i�x��n?���wy@���xZ~)��q�.������8l��ž���V��u�[	�ـ0�g~���و����~��/e��mr����Qf#�4��B����%��o�~�B"�0e݅����8[�����_|i�ǳ8ήK,��������di�BVZ���ǅ���<^@����_�o��˟�����J������$k�?�}R�?����k�{�ܫ���/��>���<w��0|�p.��\ٞ3:���������IQ�,1�I��6|�g��:7oq�t�g�ۯ�>a��O�.�ro:�?�#n������m0G;�)|����t�F�rQ�e�qp�~ ��POc�Pe�H��w��^)h�ɫ��#�h��L��+v2��7.����e��a7�yy@��q�×��|W����q7�< ��qax.�|y��'R,�SO����I���[�)��m=��P�ߕy�f�3�SYw%e�Tu���c֒u�;y[�:�|2h��oL��h�~����1@��5��G��GW�K�����-Yq��Ǣ*���+ߌ_Z����;��m�jJ9>[�X��m�ʸqD�/��k��L�_s�޲5{�|�S�W��7]zi�����H�ɭ�kQq��I�I���H�{<�Q�:�z'Yzi�da��diȌ��|���&����޷#�oz�����׌��Mm��Ѭ�����f�4bF�W��t�M���m�oG����ٻ���LY�y��w���aČ�+ ?�:N#L�����"���9�Ґ	�l�����E�h�^Y���1F�(���ӳ7x���-����{޽6{7_�:W��[��/-����9�Ґ{W�+��	���?T�*}��M�;��|����8��;����űp�W�Κ��_iVt������d]��s}U�����Q˓1WwW�3ӽ���~�˺�qc髇�}(�����1�~}���g�������PK   ^IT/�|A2  �2  /   images/c4024080-3c56-4e5e-b45c-9055d78fcf58.jpgm�ct&��6|�N���ضm���67���ƶmkc���y����ou�93�S5�L�T_ݧ�s�� (-.%  @�
�s��������������C���!�b�ѐ0PP1P�А��PаP1а	q��h��HQ��Y�9ȈA ��������h��h蘈И�@ 2&� �	� ���CC'���� C����!�"��!�| ��A���
� �_�j�\��� @�`�/�!��xQ�%��O�z �ßD���1o8��{����vz���!����k��{(l�f&ņ[h�z��?�y����`�h-x)>�Y��U&��*t�#�6���Q6N�6AC#�����7k�w"��N��w���;�{������������-�^uD���m�>]�I՛k�ljq���o��J�%���(�ޏ%則��N2��;���Vv���>��t%|��Q�~D8��V�_9F�õYΘ`K�i�~otR��_ų����K�D����1��s ��q�/�mk��%1�]�~���:s*G����P�si6�e۶|�ŗk�oTǤȯd:ФY��7I8� ��3堃,.�I�%L�R�f��\-�,��X�ݫ��[�W8�����>��$F�sv��3�����G�mr��vC|p�k���͒��9m��pv,{���t\��@�:��̜�Y$�w/0ނ���ѝ��b�Ǒ���iє^{��n��¢m��b|��`�n<��3����#��#�>���L�ڜ�[�T��H���F���wxw� �cp��Y'�Ɍ�GH�y̯��a���%�g��.�d�$5��M��;���I�+�(Ϋ�������S^��Չ�5�m��+l��:q��i�����6��	0��i+C:o����8��~1�(zuG�xSMCn�&�%��|�j-�/���Rn��Ӷ7�[uS�8'i)�ݹN4?R&�H�k���=6���ˋ����y����P%�{;9k%��|Ϥ��j��������CE�c^��Ĺ�}��S3�G������5��[":7(C��$[6��=��m���:x�n���f��3 ��1Ȗ�f�-�بw�=U�nt�e���,ʇ�d��oGs�zz�1�!$p�
��Z���X���}C�]�0�tS�-��$ͣ� ���B^vҏ�ٽ]v�e��}DWL�:uV=: 2��ݢ#^�ᤒ�1֏��5��(Z|[i�8C�0!����M�ݩv¨y���r��%x�2�q)����e�t��@���ad��)aY�F4���Tұ�,���T�2���F�ڋ�jc�%{|���!
���A��ͯ"��d3{������:��2�q�KM���$�?s�^M~�)�k��6�4����)�R��Y[���������5���eʋ�,>s1G䱩�=�BH�U��=����x? �L��RZ�*�`!�����ruX%;E5!w�}��������-�Tl!�(����I�����Q
P(W���+Va���I������ޚK��<�x_t���3DMg��?_��^7�<ˣ]&q�v�9Hx��o�q�t""^�s��l��<��~�j����_�,�򚘧?d����2u�^�� /�z4� ��_@�@����A��+h�~)��!PP��"BbF&fV6A!R%aEG��8�� Р� +q�#v,���}'���);�b�8��/��k�F���N����_G���=;����]G��tx���Ťj~�yx�{t��*Rj���b����~E[5�����u��q�S�����ɡ��(+Xc��<�+��OavAi3�������$����R���\������[����	���ցgTM��v�Ã����桙]t_q6׮#1
���9R�o��>铆�:�|��ƪ������S��9"�M�\iU�̀́�9*���:QkI~�'^0��ͼrX	�W_��d��U�P�T�~�Vr�Y�����V>>�H)�����O�oE�~�����5�$��-�/�>	�^3�����}gJ
87���heP�	��3~���G��tX$8�a��XC\�}��Bկ>�]��Ʋ6�Hت�¥N?,"(,�Ŧ|▣J+%�������:_����Wd�$`�,;U��˟)��jB���:���f���@B'1��j:���]����KK���Mn$�O3����˻���3��jt`T������>x�TD�������?�Hi2�$D�k�}���C�c��e����;MHw}����^����d��b"��'	g�Tt�ư��]��
����EhGf)��Qw�h��tlq�-�V�#�[�4	��������f�v5��ғ%�����>k�9M?m��(��/W���a�^���]\\�,%v���M�5
R�����-}�u*2�q���z�T��U����j[F�f���W�� ��n\�4t~��y>O5i���oC����n^NBx����l�a�0�
�1"�N��u�����5���ɚ��R�8��T��1׼�l����4S�?j=\�����U��:h�*Y�IhG�-UT)k�S��XoP��oP_�yu
�lu7u�*�g�1~Ѭ�F��T׾���HCW�n@��c4��P��d�s�&g�x5(V|��2�c��H��j��BY +�QM.�SV�}p9xw�.��.��T0��؂�\NgwlPs��ZCj�x���a����G�L���?��YQ�n	��T�ڤ��L<'��Jǹ�i-�V�3����@[Y�Rｪ���4*x����U�<}�����J�U}�"����+�2 �d|�r:tA�P�aܕ�u�m�����{�0ѓ���i�I�t��K�̴�M�܄�NKV�����gw{$�7�Ԧ��8���X��4��e�!���F���/Ť��8�%hT��X�1�'���b�V�\]��Ry�x�N��h��<�c���J[[/�/V�;�[HN��*�����SY��D=�/?�آ��f�l[ ��x�,n�.N�.�k�}��\�W�3�ĴS�]��0Ű�ʂJ��ڣQb� =Sr���;'��1'�<��	L�"Ŧ�g#�:&M��/]QH(	��]�7�z���_^�&w,^=v�@�`aMmo��q�766>�	VP�ꮅω�&NH/��4����K����;V�Ӌ�w���U�<��" �KN��W��*��tU.�~��̪N���Ji�2\�@B^��J1q�E�>�N�C���3��f�7W�`�I���Oy���o��j�<k��;�T��,����<��ʼ��V^v�*��^�&J4�9&	S�ȈHa0�oH���H��V�A
e��^���)-��r%4�.�R��q&2�!�&�WW�É��?�i���Zif�n��W����q�<��է��җ��~�P���E��W��J*I3������ތS ��\9�$'UG�2h�ԀMA姰Bqk"خ��V"��Ş�C�&c���8S�Z&_�L�T�T۩�K=�����ķs�:bB�-W�7��3M*��N���K�����9�4�*�3�b�� ��~P�h��Ә\�D��*l�Z��z��u��Y�O�7����}�bc�B*�j�z"���Tk�S-9�OC�a��_�U��������{3o0j�b
��f�?d�Y�eQ��D����7s��s8�k�"�B#>�+��O����&�������I�s�\X;��'44�1,�����7���|�!�y�ٶ�2��+.���r�*��jX]�v=���޳�$�~�+�/��$�!$\����U�Ig��zȷk�����v�;Sa��������s��jP�H�(���m�S�ʝ^�}��$���������R���leC�Wb�����%��\�9Ԯ��:����%���T�08�)T��Aʳ���0��Q{��2Ƈ���JB��t�F��A�tl�l�mk��ɚ�G��Q֍tlh�K���׼�OU�[V�G�r�3�T�d�&�����?��������/�E� �"^`�;UF 	����@�ö@A@�1<��x�{\���#(K��V��x����{j]�B!Y]Q�3��$n�0W���"�K�TF�;�TW�T�NmD��O}{1�X��ՃhJb��*r��+�	�F�� C ��}WuXC"_H���0��A��/�@F&!PBAE"b��@�������M̔JIZ9�Zj�Ħ�zUD_azur�VN�V��(���^.*�d��vw�U��������<F����_t1H�50D:���;��Ѫ�C�		ɓ�4� ���?� ��`(DLJ@bf!C��:BFAeǼ�+pT��#'�k�����f�0����FF�rTEL�-�ŉs�驩_55]E�R�k8i��b��5fݭ���5�7�x�u�Q,^���Η+�s4��ի<5���V��
�O�9j1�ޥ7Zj�j�`�Z�b�A�AZc���P~!��]~c�4��f;�\�.mJ/���}SP0m[�E�_�^4Ť��+d]���S�^飧N�m�f5+�i�	 �P9��f{T�eu�/���AF?�����I�¨�O�W(��������Tg��I�䰦g֪cby#��u�@����:�a2�a�<�����{9q��M�I"�9_��+�<��*�T�}�H�[�cdү9���cQ��e͌��%��
KZ�����f�jӍ���Kt�k������3��f:�׸�1�
=Wkӳ�;P����c��.��@��m}��m8�K����s�����,�[튿u�{�3A�+ҽ�]���gj�UK�_Ŷ�5 �J��j���r�GU_�t����A�)��[�eКN[��j��65��&��K��j�s�LE{4�AL�Z���v����h4T�a����uFc+�U[{L��.�R[
j9g�S�F�Z�� B��tZ��ꕜs]��.H#��෹�G�PW\�>T��p|Z�ߦ�ZiY,�A0�%�V�nM�)Y� ++h� lFul�$� k�َ�|�->�:� ��HR�&�ؼ�������<Y��
�D��R�'"��yhl��R	Vw��)ͭՀ������M���*�0���$
}}"������N����'�9����Ɨ�KEu�:�������@�N��˱ �z�и�7*������!1��4%Y�x�?W�L$D�]������e5���i�i�:"jt���}&N�0}�<��	���b`��z����lU2��Y<7��V9�{$�V��X���T�e�"�-V�E�7�ʙǒ�U���SO�hlm3�-��,���0�Ɠ�0�b��|4��]�
�j��DG�(��ўB@9���i�������*�@�����STu��1I���5�S.�����l����i /�-�p�G��R����FS�c�߫�E�K{�/���� B#�tq��
'��1��IQ��lҋ���������t�*�8���m6�u
d|wk�䘳��Mli�
��mjhH��y�,�v�	J�8� !�~�[��pq�;����H����������]+�-����iv��#����j��]�C �΂�;�"g�]HF����E�I=ʲ/F4G�N%{4�A�k��&:=� 窍
83�ׄ���m�]���'t��gB�
�6��\�������8h�RInG|<(�P��O�My�v�F���iZ,h-^�ggʘ_\�`ٶoM;�ť��3�T�����~��OѸ�J(R��Q�^�����nO����kl�2��I��J}>���W�Y�1����{\��:��O'K24(�p��CV}��1ִ��<��8l��(�u=��ٗ��P��s�i	�ؤ4���ͭ���������P3���*�}���
zgW|�������ߝO�ոK�<�	�[V	��`�0I�`v�qU�!���K7�I1^���濏~a��_@��yj���$�׍�srw�=�ڿ�tr|l��z����׻t�lC�t���}L�֒��Nt2����yo���'t���8������#���C"5��W���C��J<2����#�?1��w�ZpG��s�>�!�Qަp�lz
K�J�<��,J�8�Jf���6��U���5T��I����s�柾�U�.�y�!�Ѕ���(��� _�������˼�0pz�<qY���L�ܘ]��g2?�5b����:R�/���n^��,V߅��'/�x�ƙ� ����]��)��v%C�c}�B�������"MZ5m�<<�
����g�Cy�n��3����Zկ��'̺�q�rfm�j�i�0]�V�͋jѨv�U���q �?k�~�饘z�RCp�bE���cyr�f�\�2�od�G�(B��,�O~0GIu,�Y�x!� ��]n!�Z�'���X�mL�b��u?^s}�Դ�����2h{��B�09�r;��K�$b�ۻ�J��n��B�Z}md�&��:R6�� [�Iԇ�'��Aǌj5�O�S��ܨI�����(�P��m�b^��v,A��M`�Ⱥro9�R�xj'����[ ��9��w&�~��i�c�R	L4�.a�lt�P��L>��8z��^��!�_/��M�8?�{[[�3 ��,juy�=��D�of�}A�npDb7���Mr���� 	eg�Yܽ�da	�ޔ����L[Z������3�����K�WYXN�cn����"�\��$Fl�6��m�}�;�c��,dL�e�$n�j��T�K�L��V��D�#�����+��e�[{���/� D��g�P[��C��3�67o�k2Od��)��Kh�f[��>��K폾�����{eee�Q��D��]<���y��Ӝi�"��A
d��U�JT��Zi�)�8ЙavDX���lR��v+���B����{�y<���^R��/��,%�PJs�����(�&��Zz4x�+����Zn�E�%��3��ja�?P���6�J7�V��tƹ3���G
��G&��v|����\^;ǀ5.M�P�Eͬ ��dE��(	̹��(�4VK����%j��㚭�$��=H+S���A��-������-�S�	6�»�l���Q+�ÕqQsQ,o��/�	����7��웕=��v�!P����'ȋ(��Qh*�b�����c�#�� �ƫ���1��B��YD'�Ҡg�,��Nu��4���A��wbU�J-V�s���д�1���;;�V����:V
榉(�z�]j���Fw��Gͦ��Z�u�Q�R��<a����0T�p>�!^�\�j#��;jR��>h�W\DV����IT�q\�*	�@�Es��+�%!��<K�	��pA���z�5~!d��2��D�,�6��,���UO�	u&��Ǻ*4��W� բN���}�����|%1X�ƁA��7=&�&�[�&�4�,D�Ҧ�ь�"���;��R?�Z�k_����NnT\�Ӌ!S�o�j�{�%:թ�Lڀ�z�	�Y�4̮df�Z����I�df�d?N��7��hQ��p��z��n�F@�&��E	��G	��UfC��4�&i;9��#�xw%^�`��U:5`f�>��[�۾���Y�!"���N�q��ʰ������ҭ��J�A�W'�����L}�TB�h)���i�G�4�J�/�eq[�ǳ�����&͛������F�&�;�X�}����q�J&T(yf��DM���n��`+�7z�<M:|&Zn<�w�h���ms����؊�I.hF��p��H|o;4�ƙ��,
�]�&�4�>n�s�r�5��Hq�SQ��$&�B���f6�T���Q��7$y�N�xt$�~���J�\�����|�%�K�`��Imk~ܒM���dD�ؽ���<����Ԛ�g8��݉_�Y:�����[��g`�o�C��,�@�������s,1���MJEB~�Xh�s+�MTD�AVu�]і��f��+�-.ͩ����wD��U��q�����b"�i^�NH^�צ5�Y�^⩮o��=I1��DX:�U��Nsݷ�&���*�ς����g��%t�J֯�Qssj�UBW�����I�Y��"
�*�|�`U���T3vd1R�:�ݩ�*��(�'J��������yH̱}��Oi�'Y`%��8z�)Jy�r%��ê�حm����Ft����E�T�H��mIߺK��/3(�i,�ĉHK@���PY�/_h�Z�QiQ�ȝmg�$�E�]nIA�&�V ��a�'k�TO)x��۹�S�4�4���\$}hw��]�RQ����g�z��w�����}#,K[��Y|�T���/äW1�Vw����M�$ǣ�r5ҳ<�Q�!\���s�
�09d|�UT)3[�{�+�\?66=�������%_�d����h�n^��<�t�lA)�����V|{��щ��h��f#J1�' �wEA��l����@b�v�'����2�2��p���/��pز�y�B"T�D[Ocm�$�ߺ��\��=P�I��7�V~��eh�<͉}�`ɕ[�,!��2��o�և�	�%6�''��6^Lډ��j�COI�����.Ԅ�Q_��l?V��+` ������r$Ҹf�㓢z[�c�J�X�J�"d��*ؙv�����,��:�S���5C�����4X�B0�G<Vi$�f����I�������O������O�o�EGϬ���H����aB�D��0�+�5�b0}*�j�K��-X˅h�Z|�(z�����+�*T��J>���� ����yA �(/��������2�^]���~RX�	��0��'`�wJ@��y'���.P�3}Iq��rH�����vg>;��V0��g��J,��Yޝ�ƟC5�oW���f�T�V��眷�@����K �����5*����; CD�6�C�_��Â&u���V �g��=*~�I�S��
2��
��sXVN�}z}p ��Ɗ�f�P�ԁ.�-.��4��\?��#���17��H��߳G�����r�8�L��ی�u|����<+<�pQ,2��W�üli��d�O_Q�rj�)}�
������h5�+�L�Qi�1$0e3Vޛ����18�k�,:ؼ����kxPS�(�C�|ts�P=���Yf��ۻ#��������Z�Q�-d?��ǯ5*�j� ��;��EYp�d�d�1(,1Jk��A0YbG�*�^��T�|od�!��9���!L��_Q�n��=L�Us���
��dG��I�~H���ޜ��DgP�bi�nt���޴%l��$R�rs\�g�Qg���w����ٕp����� +Т-�`��}��A�#�~���wüS��ƙ��}��*��ЙgAYF)�߀{0��fu���%b��
�c��A�K�k�����bNͻ��ﰠ���	y�v����ݩ��R����.��t���x�W٬k�����5M��-�?�~�B��ҩU1�c�.V1؅����fhyҥ}В��EW��9�U�4*�;����=�/� �Jl���^���\m�؉����7�Ȝ�d&�X��������U
�:wq~-���������'j"�F�͏m��?��j�zf�I�[ܔ�&^��!v�tX�l����#�%y��l��D�%s����3|��6d�^{�9�a����{Y��v|B|'�\��՟q�vNio��Ӹ_��'RK#5p�0�c{'�o��Ň̛86RMy__f?�p��/�R W�FT�W���$��!
|���n���Ș[mw,K����N���c{���Z
��)�*$6Բ�)�{�c���{���3�bA������p~�-���u�,���m�j=�`���!�c��d<[�)ڜV W�h�M8I�Bu�1��4�lB����`M/���0������'��gu������� �h/
��a��]	NI���RbڀC1��g|YENYjr*s7dM88�WI�Ͻ��a����<�z���pQKG�_؀�bI��%����_5��d�L�����.ᠬ��JQ�ϡ :1�: LV@���K
e%!�M+H��U�6���u�;��.��Fs(��ī��X�'���k*V����I���w�_~���3��~����ph��	@���` �xJ���o-��$O~�/oӅ�h�����T{���O��4�0+
�:AY�]��܈�-���z�(�y�D�;p�1̾�+�F�7ƀ�B��y��T@�Cqm}��K�q㼵H��F���e�b�l��<�,XC$;��ܵr��U��yLV�B��n撷Y\�I~%�.|�i*�&�:n�dn��p GE"h�<	E��#�ь�|g�"���ޣ�' ƽݡ�xTe�0��0�>�8�{lMI$���h	��CgM���w*�$��۱^&�so.�U���8;(�ҍ
}X��/���Us�÷�S��؉��C���;MЇ��X]�	&�Ns�فY|xx��)�� _-��K^��2�gSp��j8*[(ٺX赕���"��N����>�A�kql9q�Ap����|�Jj0M�ѢF�ݮw����ÿ�S��
��RB4:�2�T�����itM���F�y���nє� y:=�e�\��Bkq�2��vҩʈSV~��=�L�O��"E�;�3�\�t�!"^��R2�w���[`ǈw8흆���;{�#u��[P/�?�l��E��E�ҳ��3��_^[&��5�m:��x�F�JE	�6n��ިT_mw3�<`:#}�p����@aV�Q>[t��SnU���Ŵ^#r�l �����F�w���Dj�W����p��S��yɚ��{�+�%#�8��B���V��o9������"������<8l�3(����nZ�%������(�X��eFۙHc�L/���RL�~O�oo�=	�~�5���<CX�D��|�А�����8ܚ����"�L:S7T~��`���Fi#b�IW_-+�Ū� �|��U��fRr�i��' v�;���B�o4	D)�Ԃ���a�U�$�o5V��RW��[�c.�h*y���Ie ��&�E�
N׹�.��c����2�O/9=3s'�Ԁ�mP)���=�ÏDcK��d��I]�)�~z�M��TRu^���<Jy!ȓV�Ga��f_W�4�=ޘՀ� ̤��Ә���m�1��9��Y��zO�Ä)\aN�;�ǉ2���t��e���J����Fk�u�0�eg��h*d.�[a�x<���IR3[����C9lW���=<�T2!T¸��y���ʵ����LD�ϛ��0u���[?U����O5@=��>V��C����<"+�r�1�;,�;�~�&8�1��a��19�R
ђ�#Sw̲��hERL( =Z��D��/��T�A�z8��; ��ȓoE���򥳜�)��5��a�(l"r	�����LhǦ�[RWSR��ux�w�)����'|��M>�E�(ܨ��!e���`:���d�]�����lca�A�2���Ze�����-b���/b��`]hؕ3��Hv�bg6�	�e[P�?�vB�?a�	ɗ2��)Х��h`���7#���GG%uV��ۅ�Q��@���U>��ޙ'�̧�F�饦���<�{�L�wYuHA��'�"�0f��P�����m����-�`ɏ���=����MѮ�=����_uU�W����:��a���萅�;����r43��=YEX�"�ؔ�%q�jh�M{��6x�ob�V,���n\<~�X��0��{���z��@���=v@瞓>7-�a�x �\�%� �$D�s_$3yt�vX]���9�X�ԏ����TV�����<4���yfm��)^�Գ��������l�4�K��D����,BL|#:8���1)�T�x��Qbn��%㞝��Z�*�%9�ݿS=z��Za�(��ߵur/"zO����䩮?؎�a�U��Z� g�ɬM�[/�h�E2�ƣ�4fL�6�[XN^'|/��`�wzmV�=�6+ւZ����F@�vW�e~��IX�,�oM�'W7i��Wq��FνA�7Vy�=�0vF�[J���s���mK\|������V����s�	YW��9��HEc��E&�k�Ka`ݸBD1�i\tIÞ~{�55n�o�#�� 3E�z踛�����<�@v���;Y�q�BF,i{���9{�	�@I��sЗj�r��LP��I��Ĥ��F���΋E�W����$
8����[�>��i�:��jS���]ͼ�8��43Nio�nZ�}�_�_��1�ܶ�?�q��^qӔ�%Ի���z?!�E@t�9��LV�J�1��uNMM�U@���JMM5���tIM�*tR�!)]��1��8��6����o�ؘ�����VV0�R��'|ͪ��ė��X�����4 �t�ڦ<D�RA=���~��`�ۦ���#���(��bY Ny���{/��LxS�7�� �"������=6�d��!{h�2��W���0	/�Sj���p�g����o'���߯��<�'��2 ��R4  %A! �H�������I` ��P�vs���.�:b���`���I� 0����dE"bA% ��1�n���<��|�Y'���Ò�!ϮcY�;pY���\�� PK   ^IT[��$P  �     jsons/user_defined.json���n�0�_��X�qȭ*����*Tǡ[;��"���]C)�Jsrvg>�׻#a�iR��k�V���IB���`6e�c���(��|��u�W���C���^Y�E-yA�h�^$jt(Ʉd��U��Rg:]�L�S�eu1iT�M�C�ep���1�^9��!�)��+���[��37�%厘~=ߵ��ֶxO���U�֣�Ė�Ŕ�[8̤7��c 3�����Ë�!漃+�咳D\SԀ�1��:t/�VKdH.��9[0�T�l�S����T��..�9�r"e��OE���/��y>l�>�%g;��w)n����6,�oPK   ^IT�<w�&  ��            ��    cirkitFile.jsonPK   ^IT/�|A2  �2  /           ��?&  images/c4024080-3c56-4e5e-b45c-9055d78fcf58.jpgPK   ^IT[��$P  �             ���X  jsons/user_defined.jsonPK      �   RZ    