PK   5tGT��P��#  ɉ    cirkitFile.json�[o$GrF��A�N2�������>y�A(��(��1�G��Ψ"�떹q0`�]����a0U_Ve��7Oǟ������w?�O_�n>I��������ۯ�7����c�����7�~���]���NO��rz�s��=�ᴯw���:U�ݩ���m�&���oo�.t���w���Ĭ:13XBW��
�+�V��Uf�B�j3�U!t������������`U���`U�5�^(��(��Z)�bi���ri����i����i����i����i����i����i���V��i����i������v��i����i����i����i����i����i����i����^;���^;���^;������Y�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"t��v�%"��v�%"��v�%"��v�%"��i����v�%"��v�%"��v�%"��v�%"��v�%BW�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y"R ��쵳��N�D���N�D���N�D���N�D�{�4KD
{�4KD
{�H|~���=���r�>?����_H������t�҅(��N�ءt�҅�`cW��C鄥]�Ʈdc��	K=���J',]��`cW��C鄥�W{6v;�NX�������ءt�҅�ecײ�C鄥݁�݁�J',����΂��O�g��G��^��B`�!��`���wH���.���O�~��;�O`>}o��6X>���c8~��`���w��������O���;�O`>}?��>X>����zx��,��|�' ��?X>��t7?�	����?
��|��8~��`��ӽ/p�`���	̧�v�������O�����'0����O`>����,��|�;~I�,��|����?X>��tG ?��|��^F8~�[V�kV��(a�Q�����O������'0��|����O`>ݳ��,��|����?X>��t�4?��|��o6~�?X>��to:?��|��z8~��`���~ p�`���	̧����;=����`�Q�����O�G����'0�������O`>����,��|�k��?X>���K
��,��|����?X>���3?��|�iO8~��`���n@p�`���	̧}���ѻ������a�Q�����O{G����'0�v�����O`>����,��|�i��_��O`>���,��|����?X>��;?�������s9�u��N��î*�rw���|����eݟ'�eNߛ/s���z���w͜��h����;3��o��9�}������\fNߟ27m�ig̻��_��79m+w�1�&'\��7f��T��������;�Z���79�(w�1�&g��7���|����*��ͱ���痧~wh�~w�㩾E����U/i��O?i��?i���>i��>i��O>i��>i���\v��/W������1�V�zi󍙷r�K�o̽��^�|c��\����o媗6�Z����r�K�o̿��^�|c�Y�z���r��or\�|c�M�]˝o̿�Yg���79_,w�1�&gz��7����������]�;�z�g̿�IO���79])w�1�&'��:�or�P�|c�MN�ɝo�����s�;9�$�KS4��r��6ĩM���*ܞ/uۖ+�3i��O?i��?i���>i��>i��O>i��>i���\v��/W������1�V\g�|c歸δ���[q�i�ٷ�:���o�u�ͷ�=c���δ���[q�i����:���o�u�]�����:��[/���[q�i����:���o�u��7�ߊ�L�o̿י6�z�g̿י6ߘ+�3m�1�V\gڭ�1�V\g�|c���δ�V�a̿�u�1t����x��t���W��-������͇�_H(���!����]�
j�"H(�+g� ��F�!����0D�P���
���ABAM"H(�0P��6W���-Xᦔ°1a�[��M)�a�b��`�R
ÚĄ�p��8���G�	��V�)�0��BL��7w�����Rև!&��X��°�1au���8���v�	��V�)�0<��8V�K��SJax~1q+)�R
V�K��SJaxv1au���8��gLV�K��SJax1au���8��gvV�+��SJax�1qk�ܢ8V�+��SJax�
1au���8���V�+��SJaxN=���x��qJ)��!&���X�����b�nr�7�:^cu�R
Û�V�k��SJ�j
c��x��qJI["aLXo�:������}�,\u�WD�������}-\�������}g-\�������}�_\�����F�������x��k�r���>�L<XŅ5ޣ���}�`&������qU0��������qU0�������qU0���ª����B+>��n�Ol�\�����]�c���y�Њ��k�[��B+>��μOl}������>��qa.��C�{|b���\hŇV�b���Ǎ�Њ��)񉭏#s�Z��[W�B+>��������/s�Zݫ�[_�B+>����'�NOĜ�����Ǘ>�̅V|hu�Ol}|�����^>����2Z��=�>���e.��C�{+}b���\hŇV�����Ǘ�Њ��u����/s�Zݳ��b��/s�Z�{�[_�B+>����'�>�̅V|hu/�Ol��Vtz]�Ǘ�>����e.��C�{�}b���\hŇV{���Ǘ�Њ��J����/s�Z���[_�B+>�ڻ�'�>�̅V|h��Kl+_�B+>��K�'�>�̅V|h�'�Ol}|����jo����2Z��5>�u�I洕�ǗU>����e.��C�=�|b���\hŇV{���Ǘ�Њ��p򉭏/s�Z�E�[_�B+>��S�%���/s�Z��[_�B+>����'�>�̅V|h�W�Ol}|����j�9����2Z���y>�u������Ǘ�>����e.��C��}b���\hŇV{2���Ǘ�Њ���􉭏/s�Z����Ǘ�Њ���􉭏/s�Z�Y�[_�B+i���D�9�u��N��î*�rw���|����eݟ��a�TY�M����M6Se��w��B��L��^ٙ*ݭ3U�Qg�,t��TY����uP�2ٻt�k���KG���0�t�i���KǄ��0Y�tg�T��,^:�2W��⥳ se�,^:q�U�\��9ֻ}�Ly�w���wG9��KQ}�o_��T6�&Ie3i�T6s&Ie3e�T63&Ie3a�T�|�,zI*�5/-��e�w�ʝ&�����;M����+w����W�4&����i2Pf�x�ʝ&�d���;M��b�ʽt�q���K���0Y�tTo���K���0Y�t�l���K����0Y�t�j���K���@w�L/���+�d��9��2L/�F��:�,^:�1W��⥓se c�d�ґ��2�Y,�8]��ٵ��eW�!*4�1��U�=_�-���T6�&Ie3i�T6s&Ie3e�T63&Ie3a�T�|�,zI*�5/-��e�w{- M����4&����d��^H�a�x{- M��Lo���0Y���&�d��Z@����kiW]&����d�[	&����d�,�^H�a�x{- M����4&����d�;b&����d�,�^H�a�x{- �u0Y���&�d��Z@�d�,��Z��Nw}�\�����ﯺ�g�k<�_�O�����G�CBaX$@� �0,8 D�P/"H(!$�E�
�B	�a�!��°p�ABaX�B� �0.h1%���\���`��R
�Ä�n��7��E�	�߂pJ)�k�V�+�RWa&��X��¸>�0q���8V���SJa\g��:^`u�R
�=Ä����R0LX/�:N)��cǱ:^bu�R
����[I�R�:^bu�R
�S%�	��%V�)�0>�b��:^bu�R
�8�	��V�)�0>#d��:^au�R
��K��[�ű:^au�R
�CZ�	��V�)�0>>f��:^au�R
�m��V�k��SJa|��0au���8�Ɨ&��&�x��5V�)�0�`��:^cu�R��uV���SJ�,c��x���%���g��z��؟PVqaݤ��
�ՃU\XC7i�G��q�`��M��Ӫ`\=XŅ5�.��N��#�`�x��Ios$����Q\�:�k�D��U\XC7ijN��q�`��M�Ӫ`\=XŅ5t�f�*WVqa�w�}����r�Z}��'�N���v��.�1^��\hŇV�5�����r�Z}g�'�>̅V|h������0Z��=>��qb.��C�{1|b���\hŇV�����Ǒ�Њ��񉭏+s�Z����`�Ǘ�Њ��U򉭏/s�Z�s�[�'bN��||Y���
_�B+>���'�>�̅V|hu/�Ol}|�����D����2Z�ս�>���e.��C�{D}b���\hŇV�����Ǘ�Њ����y1�Ǘ�Њ��=����/s�Z�C�[_�B+>���'�No+:�����J_V��2Z�ս�>���e.��C�=|b���\hŇV{%���Ǘ�Њ��|����/s�Z�]�[_�B+>�ڃ�%���/s�Z�%�[_�B+>���'�>�̅V|h���Ol}|����j���:�$s�J���*_V��2Z�՞A>���e.��C���|b���\hŇV{8���Ǘ�Њ���򉭏/s�Z����Ǘ�Њ��󉭏/s�Z�q�[_�B+>�ګ�'�>�̅V|h��Ol}|����j�<��:u�pj����j_V��2Z��^�>���e.��C�=}b���\hŇV{K���Ǘ�Њ���t�m���\hŇV{}���Ǘ�Њ��,����/s��4�׳��ۺlw���aWe�;��yw>\n�V����K�0g�,���TY�&�����;Se��v��B��L���֙*��3U:Hg�,�|��:(y��]:�5W��ߥ�Use�^:�4W���cBse�,^:�3W��L/�R�+�d��Y��2L/���*s�By��ݾQ�<��CS���O��(���I*�Y����4I*�9����2I*�����0I*L�l�$�͚��uP�2ٻ}�N�a�w�ʝ&�d���;M����+w����W�4�3Y�}�N�a�x�ʝ&�d1t�^:�8W���C�se�,^:�7W���qse�,^:v6W����]se�,^:B5W��⥃Jse�;b&��N�̕a�x��\&��N��uL/���+�d��Ɋ�2��c�x���\��,�P�.M��������e�*ܞ/uۖ�kI*�Y����4I*�9����2I*�����0I*L�l�$�͚��uP�2ٻ��&����Z@����ki2Lo���0Y���&�`&����d�,�^H�a�x{- M������.���ki2Э���ki2Lo���0Y���&�d��Z@����ki2�1���ki2Lo���0Y����:�,�^H�a�x{- M2vL�i-���_�����񩻻�z�)|������}�?��Kw��=>]���O�}���S�������e~��������r=^����������]��w��O��~#���k�uoc�*�Y"+F
�DV2�f�0��)�aXI1R�%°c�0K�a%�Ha��J���,��$#�Y"+QF
�DW��e���D�� Ԯ��8+PC(�v�0.Z9�:*@!�k�qA���R��]#�K�V��@=�k�qQ��A܏7�@=-�zj�㺲���PO�a\ٶr �� �]#�k�V��@=�k�qu�j%�zZ�Ԯ��V����%PO�a|Db� �i	�S�F�X9�zZ�Ԯ��DV��V@=�k��A����PO�a|Tf� �L�ES��V@=�k��i����PO�a|�h� �i�S�F�xZ���zZ�Ԯ�g�V���@=�k�񩯕�x
E<��i�S�F_b�r ���]C;�@=m�zj��V PO��N5�NM��qzc[(���|�nҹ��C���	��Iw2N��'0_�&��9=$~,��|�o��}6~�,��|���ߤ����e���p�&훍�/�'0_�&��9=$~,��|��tc�����|�n�q��C���	̧�)�7д�	�&�w,��.�!�ڈ�D`B�	��V:���	�&��r�Ҏ&�P�)�cH��PhB}��!�L`B�	�]n:��;�	�&�����&�Pߡ�cH��PhB}��^��}
L(4��]�cH��PhB�wA�b�?2�}JA����)0�Є�߅�!�S`B�	u�Cڧ��B�>#:��O�	�&�=Rti�
M�����>&�P���1�}
L(4�_�}
L(4��	�cH��PhB��Hǐ�)0�Є���!�v�z�SJڧ��O�	�&�=�ti�
M��w��>&�P��1�}
L(4�cH��PhB��Mǐ�)0�Є�_�aE��PhB�kOǐ�)0�Є�'��!�S`B�	��Cڧ��Bj:��N|+
�S*ڧT�O�	�&Ծti�
M�==��>&�P���1�}
L(4��R�cH��PhB�ǰ�}
L(4����cH��PhB�Cǐ�)0�Є�;��!�S`B�	��Cڧ��Bj�&:���y|�<�SjڧԴO�	�&�^Yti�
M�}���>&�P{��1�}
L(4��W�c��>&�P{��1�}
L(4����cH��P�_p�rl�ݝnO�]U���N���p��[)ʺ?OO,̜?�M�9�S0s���j��IO����^���'=H3�Oz�fΟ��̜?�ՙ�?��f����\kN6��f��(�\kN���f����\s-�f��d�\k&N�r��f����W�s���X��m�������x�/EQ�u�vEL���I�W� i�J$�_I���+�4%��[�+�(i�JJ�sZ3p튘&`���+b��5׮�i�<\�"�	X3q튘&`���L\�"�	X3q튘&`�D�qz`��5�G��
X3qz�]��5����
X3qz�[��5�G��
X3qzhY��5�Ǆ�
����8=Q+W����3�r��8=5*�>ۚ��s�r��8=)W�lV��8=D(W`%%�KS4��r��6ĹM�}nϗ�m�5��4%��$A���H���I�W2 i�J$ͷ��W
Q���:��?��f��_M����_M�f�_M���_M�f�_M0�Bk&���4k&���4k&���4k&��մk�5��j����l��5��&`��5��&`��5��&`��5��&`��5��&`�C�f�_M�f�_M�f�_M�϶f�_M�f�_M0�k&>��?>ܼN��t��.*~����M�S֛O�݄H!�O���O���O���6�9�a��*:Vt��h���E'��(tF1h�Bg:���Έ���o!�`�o@���3
�Q�Rg���(uF�3J�Q�Rg�:���ΨtF5|:���ΨtF�3*�Q�Zg�:����M�Zg�C SR��8���/����桿�M������kw<��������}���ݻ�������U����_oK��x����+�����?@�ou�˿��(���>=~w�P$~�����(֓/ק��bd�?��n~>���*��Q��p�n�}���{��(z���x���~��v���t���S��_���ͧkd�1������x�~}������^1��r�}�zw���<\����ة"���/w׻���vEq�x�7u��a��� ��q���0��� +�_�F�������ߕ�Ի�R�]�owr
��r8���fe������eNB��p��Ň�qD���9~�|�t�����D��9_h�2|�!~R+e-�?)�}R�O�P=;�>i�9e��+�A�PJ��K�b����;�"�c��68V��Kux�R9��^��Ørx�c��Hю����F�}p��W�R���~�L�M�,���o|�y�S�s�v�o�S�O��c]���[�-$����7��1�c[��G�0�5ML3la�4IN�|f������]����r��������#��"�2Yaq�q�7
a9T=�P�}]�-��C��}Q�N�S���m�;�S���CQ�˺��0�/� ����������6dC�Lۼ��1�_���������yN��e��Y��������y�����������y!�� U`WW�����n�T��?<u��7M?�����v1{���%Hu�4�*Ҙ���G��/��C,��KMy[�á����79�`����[@�8�>�}	��W_���#M�- ��G�4R�T�oI7�`i:nif�<�xi��y���摦��f�"=_K�޿C��`if�<���y���_�����x~7p����y�+��y���������M�/��/I7��<�t����y�j�Q��_͙摦��f�#��w�/�0/ף�摦��f�#�weE�R����H�qH3�H������x_�Q�x�/��sY}l�mS8����.�/�iύ��iޅ�?ě���շeq,�oo��x�p��}��A?8i���>dȦJ�9G����sӇߏ&^T�g�~<7y�}o����o>���콢��������FE�����#�w�Wj ���^>�������0�16G3553l��0~1�o>��y��,���g�~n ��փ33n6K��f������{�*�����~~�,�t�<�̸y�x�Z�"���t�,�t�<�̸y�x�ʲj�~���%z��<�����V��x�{P��f�����f����0��Y/����Y�׏�9�|>��tߖ/�z)���fy���f�����xiٗ�|3���f���͍��+�7R�M-a�F̌����7Ϸ/�}�^!���x��UQ�2p�y+�O^�>\�[��c�Q������jx��T�k_�k��]�?�/�ׯ��������}?�?���������������^��]����/Ã��PK   5tGT��P��#  ɉ            ��    cirkitFile.jsonPK      =   �#    