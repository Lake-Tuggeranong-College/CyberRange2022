PK   �ZIT�� ''  I�    cirkitFile.json�o��8�ƿ������?������on7��I ȶ<1���s�'3�ݏ%��nS���S��2��L�|��R�Ģ���ű��{l6�c��������=�w�O�q��}�Ss���lN���c�����+�wv��s���]�]\���W�Y/��t�fźXe늖Y]��)�fY���4fq�����+�X�4$f�*�Ɗ�
���R�b��iJ1�T�4��A�`���A�`�Z� U0�J� Up1J(��*屒��R,�(��R,�(�S,�(�!S,�(�AS,�(�aS,�(�S,�(�S,��V��)�p��)�p���<vZy�K8
y�K8
y�K8
y�K8
y�K8
y�K8
y�K��P;��B;��B;�����cg.��b	G!��b	G!��b	G!��b	G!��b	G!��b	���)�p��)�p��)�p��)�p�INy�,�S,�(�S,�(�S,�(�S,�(�S,a�R;��B;��B;��B;��B;����H;Ky�K8
y�K8
y�K8
y�K����N�����N�����NO���Kw̎��!z�C�������]�'��c��P�|��������c�xr~Im]�u�ޭWYa�<k�z�mV�]W���nï�`(�Of� �;���t��X�Y��t��3M��]�����t.��ڮ��JGX:7��ڮ��JGX:7R�ڮ��JGX:�,��[bm�#,�ij��j��t��}�Pӊ���Ya���JGX:^�X�3,��x%�~�����s''�N�|�㵫`��3,��x�-�~�,�G`>^/�8S����W:���V�|��5�`��3,��xu9�~��G`>^�8�����W�'������|�l?p���#0� ��v�z�Xp�a�����|�sl?p���#0���`��ǻ����X>��>'�������|�Cl?p���#0�-��`��ǻ��<�����|��l?p���#0�D��`���{(��C��B/��98�������|�ol?p���#0���`���{����X>��.g�������|�?l?p���#0�,�گ �X>��x�������|��l?p���#0�! ��`�����C�Ao�8�(�����|\�l?p���#0�� ��`��ǕB���X>�q��������|\�k��`���ue���X>�qE�������|\�l?p������u�a��]]v��PU:1�e�]Q�ޮ�S������ԥ�.X>�q�%��Л�ѻ���K	N]Jp���}�W���h��+e�M�z�|��_`���,���:�~��G`>����_�z�|��p`���,�����~��G3|��Bn���u�-!����njb�ۂ���o+�&v�-1����6hb�ۢ���o�q�����H2 ~["'����_�����HP��ߟp&�(7V	����P��_�u�K�/�Byq���ra$���J�/���QQ������t�)L���2[�����]��8�Q�.��ڮ�&�Q��w?�{��Gu�����[�=|磺�o|Tw�}������6R���w\ij��yG������S/����&�zq���7�ԋ�/�{B��x������S/�����O=�8���B���K�/�?�ؼ��B��K�/�?�x���B��dK�/�?����B��K�/�	��;�+�����ñR���;�*u�,�?����B��^J�/M=���S��?�d�z[�*���6+j�V]��w��m�e]�YgT��ݏ���Q���>�{��Gu������]x��a'�{8�Ĺ���~7�u��z�D��_�{Yg\��Md�q���7�u����=��Md�q���7�u����D��_�Yg܃K�Yg\�W�Yg\��Md�q���7�u����D��_�Yg\��O�Yg\��Md�q���7�u����7�u����D��_�z�o"��* [up�kA�BR�*fD�ɩO���������l�����U.��Xw�6�����J������2H���$dx�C2<�!	������a�@B���0D !óX"���'�@!�qa�	�QJ��1�b7��7J���� &X�&X G)�~�����(%�O��`q���8J���� &��7 ��q��(%�O؃�`q���8J��/@L�8naq�d�  &X��8�R2��P:��9,���L�B	Ą�I�M���x��(%ӿL1��x��(%ӿ�1��x��(%ӿ�1��x��(%ӿD1��x��(%ӿ�1���q��8^��8J��/�AL�8^��8J��/�AL�8^��8J��@�~`q���q���8��`q���q���b��po7q�7aq���q���>��`q���q�3�1��x��(%.�c���
�CJ�ŵnk��U��XU���S���*��4�5��@�j��
�ink��U�v�`%V��V�����J*�.�R��m�j�4XI�Ս�T�z[�cVRauc��V��X@��TXMs[��
��+���涖5\hWV�~e��,���q���m�k�4XI����$:�
-����f�*e]Ji�N�E:��d^*��C�k�ul��}�В-��ױ�N�BK:���_Ƕ:Y�
-�����db*��C�{1tl����В-�)ѱ�NF�BK:��7FǶ:Y�
-����:y�
-���^%���e*��C�{�tl��FL镘N^fu�2����В-�ӱ�N^�BK:���OǶ:y�
-���D���e*��C�{+ul����В-�ձ�N^�BK:���UǶ:y�
-���]��I:y�
-����c���e*��C�{�ul����В-�ױ��jE��:yY����:y�
-����|���e*��C�5tl����В-�Jб�N^�BK:�\�AǶ:y�
-��r�
���e*��C�58Tl[��e*��C˵Dtl����В-�Dѱ�N^�BK:�\�EǶ:y�
-��r��*�$S�J���:yY����В-�ұ�N^�BK:�\�HǶ:y�
-��r'���e*��C˵�tl����В-��R�m����В-�ӱ�N^�BK:�\�LǶ:y�
-�К7�!m�����������}ҥN^V��e*��C˵�tl�T�C�̇N^v{R��,Ҷ>-���
-�2Ա�N^�BK:�\�QǶ:y�
-��rmI���e*��C�52Ul[��e*��C˵>ul����В-�,ձ�N^�BKq��GD*ݦ4Q	T�MT	��NT	T�NT	��NT	T�NT	ԣNT	T�NT	�|N�:���K�TK��O�Se0�;��g'�2`�*����1��2/ƙ*��� :�2U�CgA��`�8t��UfS�|W�e������]��l��Ԯ˭��+��'w�ʬ�D��:M�ʬ�D�̺L�ʬ�D��:L�
�_f�^��l̋�:��b�7t\{��C����`<x��'����'w�Ƌ��q2�����'w�Ƌ��q2/=�C���`�8t�p�ƋCG���`�8t n�ƋC�Φ�`�8t�k�ƋCG���`�8tPi�hD����	��2/���*����i��YƋCg>��`�8t�b�(��xq���T�Y/&c���VY�m�YQ�Pu���
��l˺����Tf�&Je�i�Tf}&Je�e�Tf=&Je�a�T0�2��Tfc^�ׁ���sq2������x��\@�Ƈ���d0^<?'��/�����x��\@�Ƌ���d0^<?���x��\@�h(������8�����`�x~. N���sq2/������1^<?'������8����e/�����x��\@�(��x��\@��]]v��PUfŚ�슲�vm��j��^�����(��vO���R���$�[/Ӝ�ө=u���W�����S>vϧc��/��y���-!	���"���c D !�O�@�@B��&���L?�!	�~�
B2�T�$d�i5H�St���ڸ����(%3�Db�`��`��d�9R,~,����0{�a��p�q���1L�8naq�d�on����⸅�q��&�1L�8naq�d�W&X��8�R2��,�[XG)��5&����QJfx��a�ͤ�R`q<��q��ޓa�`q<��q����a�`q<��q���-b�`q���q���zb�`q���q����b�ps�IqX/`q�d���&X/`q�d��&X/`q�d�W��W?�8^��8J��0L�8^��8J��0L����כ�8^��8J�;:0L�8^��8J�����`q���q���1��x��!��Rn^�@��Pq�J*���j�L ZhWVRa5�W"�
��+����+ێV�U��TX]ޥbW�b;������A*v���C,��J*�n��bW�R;����j�L;ZhWVRa5�W��
��+����+ώV�U��TXyM�Nb��q�В-�mֱ�R֥�v��]��x�N�BK:���\Ƕ:ٗ
-���y��d`*��C�k�ul����В-�aб�N&�BK:��CǶ:٘
-�����dd*��C�{ctl����В-���y�����В-�Uұ�N^�BK:���JǶJoĔ^���eV'/�:y�
-���8���e*��C�{�tl����В-�IԱ�N^�BK:���RǶ:y�
-���Q���e*��C�{]ul����В-���Y�����В-�=ֱ�N^�BK:���ZǶ:y�
-���^p�*�VTZ�����:yY����В-��ױ�N^�BK:�\c@Ƕ:y�
-��r����e*��C�5tl����В-׮б�N^�BK:�\�CŶ�N^�BK:�\KDǶ:y�
-��rM���e*��C˵]tl����В-רѱ��N2��d:yY���:y�
-��r� ���e*��C˵�tl����В-�pұ�N^�BK:�\�JǶ:y�
-��rM-ۖ:y�
-��rm0���e*��C�5�tl����В-�jӱ�N^�BK:�\sNǶ:y�
-��r�<�*U�P*󡓗�:yY����В-�2Ա�N^�BK:�\�QǶ:y�
-��rmI���e*��C�52Ul[��e*��C˵>ul����В-�,ձ�N^�BKq�ף���u���z�^e���5�M�Ymw]M6/�M��D�@m�D�@5�D�@�D�@��D�@��D�@u�D�@=�D�@�D�@��T�9/�{C����`�7t�j�ƃC���`|8tLh�ƋC�q�ʀb0ƋC�T��`�8td�ƋC'.^e6��wU[f��8�|�e��vYK��Zk���rG��zM�ʬ�D���L�ʬ�D��zL�ʬ�D�`�e6�E��Ƽ8�9/�{��q2��r��`<x��'����'w�Ƌ��q2�����'w�Ƌ��q2/=�C���`�8t�p�ƋCG���`�8t n�ƋC�Φ�`�8t�k�ƋCG���`�8tPi�hD����	��2/���*����i��YƋCg>��`�8t�b�(��xq���T�Y/&c���VY�m�YQ�Pu���
��l˺����Tf�&Je�i�Tf}&Je�e�Tf=&Je�a�T0�2��Tfc^�ׁ���sq2������x��\@�Ƈ���d0^<?'��/�����x��\@�Ƌ���d0^<?���x��\@�h(������8�����`�x~. N���sq2/������1^<?'������8����e/�����x��\@�(��x��\@��]]v��PUfŚ�슲�vm��j���'�Q*��;J����v���۩��f��mqOw�/�c��|~h7ݶ�?6��;.�߿���4�k���7��?�	P��fa| %�+D$���$($D��nP�~����Ǐ>v�~u�>nǜ�����x�G���{���Ŀ�Dh7������=n������Ԟ:�/�}����th�������/[�v�>���K��)ּ�M� ��韂B
��韢B
���҅b	�O�)����R�%L�*@H!�0��!�X���"�b	ӿ�R�%��*D��>� T�a��9R@%@�k��}��G	H�fx�%� �RS��ީI9 ���\�o����(b@
��O�fx1)� �S��r3��r ��S��^�J9 ���\�����$ ��x*�0�j)"�G���x��\��إ�x��\�o���x��\����xZ �\�+��xZ �\�k-��9SĤ) ��x*�0�r) ��x*�0Â) ��x*�0Ò��> ���x*�0â) ���x*�0ò!)�-�5 ���x*�0�.() ���x*��R� @<� �T��%�xZ⩯�^��+����
���uK�s�&�5�W	�1'���|��]�� �����4�I8=���|�s��~�1�ϋ�#0�n��� ��X>�a�~�q �ϋ�#0�i���8=���|�3�W�����[��/E�M���ӫ�/��X>��*F�x���		M�+0�6�'%���:/!tb&$4!�|E����		Mȫv�6D'(`BB�c��I
��Є�ZmCt�&$4!��F����		Mȫ��6D',`BB�
{��Y
��Є�; =o��S���&�h��0!�	yWچ�(�7(�<Ţ���S���&��0h��0!�	y'چ�<LHhBޅ��!:O��wP�m��S���&��_h��0!�	y�چ�<LHhB�u�^��S���&��h��0!�	y�#چ�<LHhBީ��!|�|�:O��yJ��S���&��h��0!�	yw/چ�<LHhBޙ��!:O��wU�m��S���&��h��0!�	y7;؆:O��w�m��S���&�*h��0!�	�چ�<LHhB�ހ�!|c
|g
:O)�yJ��S���&�h��0!�	��چ�<LHhB�V��!:O��+��m��S���&�*1`��<LHhB�p��!:O����m��S���&4o������	�o�폢#~�Hڤ�LHhB.���!|O=|S=:m�=G	*���Gx�M�q������ŀ		M�5��6Dg1`BBr}3��Y��Є\�l�
�ŀ		M�u��6Dg1`BBrM<��Y���h��#��(���#L���eM���SM���AM���/M���M���M����L���?�-$z��#���C�#ӦJX��I]�?�,U@��)a�R����JNi��J��N�ШT�'��4]6��wU[f��8�|�e��H�v]n��]�M=>��OxAT�	'��?�Q�'\ ���D��p�����?���Oġ8�;���NS�>�)�* �©'b������qRO�z"�	�c�����qRO�z"�	H=Q�D�OL�z��_����S�R���c�* �D��T�'�g��
H=�?-U@��yd�������R�����* �D�x��q����R�����* NV���V�*0�d�z[�*���6+j��V]����6۲��|5���D��p���>����Ox@T�	��/���(��D���J=p*_����T�' �©|5N@�S�j������8q,�z�T�' �ĩ|5N@�S�j�����ոg�����8�cY�S�j������8�'N�qRO��W���8���	�G�RO��W���8���	H=q*_�gK=q*_��z�T�' NV��8���K��e��UeV�9U�+��۵���rۧ�S��F�z���������*��6�C����_1�����:����Ge>^�R�+����[�Wܦo�-���%nLܚ�9q{��=,���6����r�=,�p���#D�&�P��p�=r�s����9�ȹG�=r�s��{ܣ��(�O�=
�Qp��{ܣ�%�(�G�=J�Q��{�ܣ������#���/�[�}tߺ����؝��ָN�[��}���7���^�,(��HD'�8�K��� ]d �����r	���='�OWH�O��Ս����S�Ю����ߍ�t�?����D�%{�d�K��R�_*Η��e��м:�|��;4���,�T.�n���ܹ�˛�nw�[� �b��kO��������sw<��)���G�?�[�S>���ǟ��_����������+/���ǽC[��=}:|���:����}x��ŧ�����~�н�������ع(xr�Ά���ϻvsz>vǩ�����_�����?�鯏�g��>���a�o���?8��Ϭ]�[-��V���-ͻ���j�S;#3�_��.�v�n����l�S��U��hm��v�Z�?V����>n.}"�Xw������v@[<v?�쏛��|_�gD�w�o����x���]����x�R,�+�)���J5�ɋ��,{�UN�ˏV���印5}c7dxi�`��Js�Q޷*��ʾM�\]�T}��|���(�|�_.����J�S��.�g������o<�\�C[�#�o�ܰ��|�/&	\e�@�W�o1r�_��@����h�;i����#?�ߏ�O?�����߻���աw�uA\���s¼�zDtW�{��,��p�ʫ��E�^��l��y���������7yY��m �J�b`����ʗ������P�i�W_|�����OƻQ����^���aT��Li�߂s���݇�c���k.�#b����_]��`f�:�ty�M�����˜����b���,lS �\��8y6�\`�-/1�u6+;4��ˇ�/�H�] }��8���T��^���H~� �H�q��IC�%r�8�a�o@i8�4<�(�n�ӿ0�� �4E:?K�\� �\Ei7�4�p���k@�/;Oᛆ�㝖�vWv��8��.�>�p��>d}�_�n��8��.�4�p�����j�\G���F�#����sy�\G���F�#�2�_�|qA�/�#��H#}$��_A��D8_�������7���2��ji_���������T���r���[��\Qf�.�mN]�[yyp��s�0p�C?�&�ۜ`����ma��H^rt,����J�go������V�^c��v����S�M�_;�]z��2ܴ��@e��\W�7n�/󐄭x�_UUq�^�A+��*��V��c���h�q�z0��b�
2r�-���c��8E�߷�Y�wt��[
��-�H�q
j.�:�t�Wc��r���k2N�#̪�M=|��J2v�-�H�[��&�$<���2?��}�c�ޒ���%k2N��ɪ4�9���d��[���$cMFI�a�k�\�[��^zC2��d��8	
+���x��OF/�%iqK2�d��ǂ.�_&z_ݝ�KoIFZܒ�5'�!`Y���zŕd��[���$cM�I�u�|~-��`]"os���W�����O������>�����YY�e�K7�*���ƍl/c�~�rP�ʶE�e�zg�U��fy�u��UfY���o@�N:b@����
�	?�ݎ�Ηngb�G��������=�tp�\������*���(�'�U����~{��~���?�����-Wŵ�o�=+�k_�ͧn���wo?������/���������9����aq�a��~��Ç���?�������������պ�툖��}/}l��eu�������<�؞>��_?|��������~꿵O������7/s��|����mV�;[����6���_Z�L���>,�9�|�e��c�e�eo�_��̢�l7��^�_���f�����x�M�</��� �=7�c��'��=c���/��H*F��0���w�����:IϷ��JXש������t�\�����]�Q�ZE?�ȥK�SL=��׌��`���}xN� ��V�
<�j�=�BO�7�f��yO��!?~�_PK   �ZIT�� ''  I�            ��    cirkitFile.jsonPK      =   T'    